.SUBCKT AN2D2 A1 A2 Z VDD VSS
MM9 net14 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net26 A1 net14 VSS nch_mac l=30.0n w=0.14u
MM5 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net26 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM7 net26 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM4 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AN3D2 A1 A2 A3 Z VDD VSS
MM13 net028 A2 net024 VSS nch_mac l=30.0n w=0.14u
MM14 net26 A1 net028 VSS nch_mac l=30.0n w=0.14u
MM12 net024 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM5 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM10 net26 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM4 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM15 net26 A3 VDD VDD pch_mac l=30.0n w=0.17u
MM11 net26 A1 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT AN4D2 A1 A2 A3 A4 Z VDD VSS
MM5 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM22 net26 A1 net030 VSS nch_mac l=30.0n w=0.14u
MM20 net034 A3 net038 VSS nch_mac l=30.0n w=0.14u
MM19 net030 A2 net034 VSS nch_mac l=30.0n w=140.0n
MM21 net038 A4 VSS VSS nch_mac l=30.0n w=0.14u
MM23 net26 A4 VDD VDD pch_mac l=30.0n w=0.17u
MM4 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net26 A3 VDD VDD pch_mac l=30.0n w=0.17u
MM17 net26 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM18 net26 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT AO211D2 A1 A2 B C Z VDD VSS
MM5 Z net44 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net44 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net44 C VSS VSS nch_mac l=30.0n w=0.14u
MM3 net44 B VSS VSS nch_mac l=30.0n w=0.14u
MM8 net44 A1 net24 VSS nch_mac l=30.0n w=0.14u
MM9 net24 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM4 Z net44 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net44 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 net39 C VDD VDD pch_mac l=30.0n w=0.17u
MM2 net47 B net39 VDD pch_mac l=30.0n w=0.17u
MM6 net44 A1 net47 VDD pch_mac l=30.0n w=170.0n
MM7 net44 A2 net47 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT AO21D2 A1 A2 B Z VDD VSS
MM2 net7 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM1 net11 A1 net7 VSS nch_mac l=30.0n w=0.14u
MM0 net11 B VSS VSS nch_mac l=30.0n w=0.14u
MM5 Z net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net34 B VDD VDD pch_mac l=30.0n w=0.17u
MM6 net11 A2 net34 VDD pch_mac l=30.0n w=170.0n
MM3 net11 A1 net34 VDD pch_mac l=30.0n w=0.17u
MM4 Z net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net11 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AO22D2 A1 A2 B1 B2 Z VDD VSS
MM9 net12 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net16 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM7 net24 B1 net16 VSS nch_mac l=30.0n w=0.14u
MM6 net24 A1 net12 VSS nch_mac l=30.0n w=0.14u
MM5 Z net24 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net24 VSS VSS nch_mac l=30.0n w=0.14u 
MM3 net24 A2 net39 VDD pch_mac l=30.0n w=0.17u
MM2 net24 A1 net39 VDD pch_mac l=30.0n w=0.17u
MM1 net39 B2 VDD VDD pch_mac l=30.0n w=0.17u
MM0 net39 B1 VDD VDD pch_mac l=30.0n w=170.0n
MM4 Z net24 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net24 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI211D2 A1 A2 B C ZN VDD VSS
MM10 ZN A1 net033 VSS nch_mac l=30.0n w=0.14u
MM11 net033 A2 VSS VSS nch_mac l=30.0n w=140.0n
MM0 ZN C VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 ZN C VSS VSS nch_mac l=30.0n w=0.14u 
MM3 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM8 ZN A1 net24 VSS nch_mac l=30.0n w=0.14u
MM9 net24 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM5 net47 B net047 VDD pch_mac l=30.0n w=0.17u
MM4 net047 C VDD VDD pch_mac l=30.0n w=0.17u
MM1 net39 C VDD VDD pch_mac l=30.0n w=0.17u
MM2 net47 B net39 VDD pch_mac l=30.0n w=0.17u
MM6 ZN A1 net47 VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN A1 net47 VDD pch_mac l=30.0n w=0.17u 
MM7 ZN A2 net47 VDD pch_mac l=30.0n w=0.17u 
MM7_2 ZN A2 net47 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI211OPTREPBD2 A1 A2 B C ZN VDD VSS
MP11_1 net051 A1 VDD VDD pch_mac l=30n w=170.0n
MP11_2 net051 A1 VDD VDD pch_mac l=30n w=170.0n
MP11_3 net051 A1 VDD VDD pch_mac l=30n w=170.0n
MP11_4 net051 A1 VDD VDD pch_mac l=30n w=170.0n
MP31_1 ZN B net037 VDD pch_mac l=30n w=170.0n
MP31_2 ZN B net037 VDD pch_mac l=30n w=170.0n
MP21_1 net037 C net051 VDD pch_mac l=30n w=170.0n
MP21_2 net037 C net051 VDD pch_mac l=30n w=170.0n
MP21_3 net037 C net051 VDD pch_mac l=30n w=170.0n
MP12_1 net051 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_2 net051 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_3 net051 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_4 net051 A2 VDD VDD pch_mac l=30n w=170.0n
MN12_1 ZN B VSS VSS nch_mac l=30n w=140.0n
MN12_2 ZN B VSS VSS nch_mac l=30n w=140.0n
MN11_1 ZN A1 net022 VSS nch_mac l=30n w=140.0n
MN11_2 ZN A1 net022 VSS nch_mac l=30n w=140.0n
MN21_1 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_2 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_3 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_4 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN13_1 ZN C VSS VSS nch_mac l=30n w=140.0n
MN13_2 ZN C VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT AOI21D2 A1 A2 B ZN VDD VSS
MM5 ZN A1 net027 VSS nch_mac l=30.0n w=0.14u
MM4 net027 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM2 net7 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM1 ZN A1 net7 VSS nch_mac l=30.0n w=0.14u
MM0 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net30 B VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 net30 B VDD VDD pch_mac l=30.0n w=0.17u 
MM6 ZN A2 net30 VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN A2 net30 VDD pch_mac l=30.0n w=0.17u 
MM3 ZN A1 net30 VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN A1 net30 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI21OPTREPBD2 A1 A2 B ZN VDD VSS
MP11_1 net037 A1 VDD VDD pch_mac l=30n w=170.0n
MP11_2 net037 A1 VDD VDD pch_mac l=30n w=170.0n
MP11_3 net037 A1 VDD VDD pch_mac l=30n w=170.0n
MP11_4 net037 A1 VDD VDD pch_mac l=30n w=170.0n
MP31_1 ZN B net037 VDD pch_mac l=30n w=170.0n
MP31_2 ZN B net037 VDD pch_mac l=30n w=170.0n
MP12_1 net037 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_2 net037 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_3 net037 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_4 net037 A2 VDD VDD pch_mac l=30n w=170.0n
MN12_1 ZN B VSS VSS nch_mac l=30n w=140.0n
MN12_2 ZN B VSS VSS nch_mac l=30n w=140.0n
MN11_1 ZN A1 net022 VSS nch_mac l=30n w=140.0n
MN11_2 ZN A1 net022 VSS nch_mac l=30n w=140.0n
MN21_1 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_2 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_3 net022 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_4 net022 A2 VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT AOI221D2 A1 A2 B1 B2 C ZN VDD VSS
MM11 ZN A1 net038 VSS nch_mac l=30.0n w=140.0n
MM12 net038 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM13 net034 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM14 ZN B1 net034 VSS nch_mac l=30.0n w=0.14u
MM5 ZN C VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 ZN C VSS VSS nch_mac l=30.0n w=0.14u 
MM1 net17 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM0 ZN B1 net17 VSS nch_mac l=30.0n w=0.14u
MM8 ZN A1 net29 VSS nch_mac l=30.0n w=0.14u
MM9 net29 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM4 net36 C VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 net36 C VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net56 B2 net36 VDD pch_mac l=30.0n w=0.17u 
MM3_2 net56 B2 net36 VDD pch_mac l=30.0n w=0.17u 
MM2 net56 B1 net36 VDD pch_mac l=30.0n w=0.17u 
MM2_2 net56 B1 net36 VDD pch_mac l=30.0n w=0.17u 
MM6 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM7 ZN A2 net56 VDD pch_mac l=30.0n w=0.17u 
MM7_2 ZN A2 net56 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI222D2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM14 ZN B1 net075 VSS nch_mac l=30.0n w=0.14u
MM15 net075 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM16 ZN C1 net067 VSS nch_mac l=30.0n w=0.14u
MM17 net067 C2 VSS VSS nch_mac l=30.0n w=0.14u
MM18 net063 A2 VSS VSS nch_mac l=30.0n w=140.0n
MM19 ZN A1 net063 VSS nch_mac l=30.0n w=140.0n
MM12 ZN C1 net38 VSS nch_mac l=30.0n w=0.14u
MM13 net38 C2 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net50 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 ZN A1 net50 VSS nch_mac l=30.0n w=0.14u
MM0 ZN B1 net62 VSS nch_mac l=30.0n w=0.14u
MM1 net62 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM4 net37 C1 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 net37 C1 VDD VDD pch_mac l=30.0n w=0.17u 
MM5 net37 C2 VDD VDD pch_mac l=30.0n w=0.17u 
MM5_2 net37 C2 VDD VDD pch_mac l=30.0n w=0.17u 
MM7 ZN A2 net25 VDD pch_mac l=30.0n w=0.17u 
MM7_2 ZN A2 net25 VDD pch_mac l=30.0n w=0.17u 
MM6 ZN A1 net25 VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN A1 net25 VDD pch_mac l=30.0n w=0.17u 
MM2 net25 B1 net37 VDD pch_mac l=30.0n w=0.17u 
MM2_2 net25 B1 net37 VDD pch_mac l=30.0n w=0.17u 
MM3 net25 B2 net37 VDD pch_mac l=30.0n w=0.17u 
MM3_2 net25 B2 net37 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI22D2 A1 A2 B1 B2 ZN VDD VSS
MM10 net043 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM11 ZN A1 net043 VSS nch_mac l=30.0n w=140.0n
MM12 net035 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM13 ZN B1 net035 VSS nch_mac l=30.0n w=0.14u
MM9 net12 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net16 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM7 ZN B1 net16 VSS nch_mac l=30.0n w=0.14u
MM6 ZN A1 net12 VSS nch_mac l=30.0n w=0.14u
MM3 ZN A2 net39 VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN A2 net39 VDD pch_mac l=30.0n w=0.17u 
MM2 ZN A1 net39 VDD pch_mac l=30.0n w=0.17u 
MM2_2 ZN A1 net39 VDD pch_mac l=30.0n w=0.17u 
MM1 net39 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 net39 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM0 net39 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 net39 B1 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI31D2 A1 A2 A3 B ZN VDD VSS
MM2 net035 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM3 net031 A2 net035 VSS nch_mac l=30.0n w=0.14u
MM4 ZN A1 net031 VSS nch_mac l=30.0n w=0.14u
MM0 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM12 net16 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM13 net20 A2 net16 VSS nch_mac l=30.0n w=0.14u
MM14 ZN A1 net20 VSS nch_mac l=30.0n w=0.14u
MM1 net47 B VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 net47 B VDD VDD pch_mac l=30.0n w=0.17u 
MM10 ZN A2 net47 VDD pch_mac l=30.0n w=0.17u 
MM10_2 ZN A2 net47 VDD pch_mac l=30.0n w=0.17u 
MM11 ZN A1 net47 VDD pch_mac l=30.0n w=0.17u 
MM11_2 ZN A1 net47 VDD pch_mac l=30.0n w=0.17u 
MM15 ZN A3 net47 VDD pch_mac l=30.0n w=0.17u 
MM15_2 ZN A3 net47 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI32D2 A1 A2 A3 B1 B2 ZN VDD VSS
MM0 net046 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM1 net042 A2 net046 VSS nch_mac l=30.0n w=0.14u
MM2 ZN A1 net042 VSS nch_mac l=30.0n w=0.14u
MM3 ZN B1 net030 VSS nch_mac l=30.0n w=0.14u
MM4 net030 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 ZN B1 net17 VSS nch_mac l=30.0n w=0.14u
MM9 net17 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM12 net21 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM13 net25 A2 net21 VSS nch_mac l=30.0n w=0.14u
MM14 ZN A1 net25 VSS nch_mac l=30.0n w=0.14u
MM6 net56 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 net56 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM7 net56 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 net56 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 ZN A2 net56 VDD pch_mac l=30.0n w=0.17u 
MM10_2 ZN A2 net56 VDD pch_mac l=30.0n w=0.17u 
MM11 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM11_2 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM15 ZN A3 net56 VDD pch_mac l=30.0n w=0.17u 
MM15_2 ZN A3 net56 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT AOI33D2 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM8 ZN A1 net050 VSS nch_mac l=30.0n w=0.14u
MM9 net042 B2 net038 VSS nch_mac l=30.0n w=0.14u
MM16 net038 B3 VSS VSS nch_mac l=30.0n w=0.14u
MM17 ZN B1 net042 VSS nch_mac l=30.0n w=0.14u
MM1 net035 B2 net039 VSS nch_mac l=30.0n w=0.14u
MM4 net054 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM0 net039 B3 VSS VSS nch_mac l=30.0n w=0.14u
MM2 ZN B1 net035 VSS nch_mac l=30.0n w=0.14u
MM5 net050 A2 net054 VSS nch_mac l=30.0n w=0.14u
MM12 net21 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM13 net25 A2 net21 VSS nch_mac l=30.0n w=0.14u
MM14 ZN A1 net25 VSS nch_mac l=30.0n w=0.14u
MM3 net56 B3 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 net56 B3 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 net56 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 net56 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM7 net56 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 net56 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 ZN A2 net56 VDD pch_mac l=30.0n w=0.17u 
MM10_2 ZN A2 net56 VDD pch_mac l=30.0n w=0.17u 
MM11 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM11_2 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM15 ZN A3 net56 VDD pch_mac l=30.0n w=0.17u 
MM15_2 ZN A3 net56 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT BUFFD2 I Z VDD VSS
MM0 Z net9 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net9 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net9 I VSS VSS nch_mac l=30.0n w=0.14u
MM1 Z net9 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net9 VDD VDD pch_mac l=30.0n w=0.17u 
MM4 net9 I VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT CKAN2D2 A1 A2 Z VDD VSS
MXM1 _SP_11 A1 _SP_19 VSS nch_mac w=0.275u l=0.03u
MXM2 VSS A2 _SP_11 VSS nch_mac w=0.275u l=0.03u
MXM3 Z _SP_19 VSS VSS nch_mac w=0.14u l=0.03u 
MXM3_2 Z _SP_19 VSS VSS nch_mac w=0.14u l=0.03u 
MXM5 _SP_19 A1 VDD VDD pch_mac w=0.18u l=0.03u
MXM6 VDD A2 _SP_19 VDD pch_mac w=0.18u l=0.03u
MXM7 Z _SP_19 VDD VDD pch_mac w=0.17u l=0.03u 
MXM7_2 Z _SP_19 VDD VDD pch_mac w=0.17u l=0.03u 
.ENDS
.SUBCKT CKBD2 I Z VDD VSS
MM0 Z net9 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net9 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net9 I VSS VSS nch_mac l=30.0n w=0.22u
MM1 Z net9 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net9 VDD VDD pch_mac l=30.0n w=0.17u 
MM4 net9 I VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT CKLHQD2 Q TE CPN E VDD VSS
MM30 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM28 qf_x clkb net0190 VSS nch_mac l=30.0n w=0.14u
MM22 net11 CPN VSS VSS nch_mac l=30.0n w=0.155u
MM21 net11 net51 VSS VSS nch_mac l=30.0n w=0.155u
MM18 Q net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM18_2 Q net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM14 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM11 clkb CPN VSS VSS nch_mac l=30.0n w=0.14u
MM31 net51 qf VSS VSS nch_mac l=30.0n w=0.14u
MM29 net0190 qf VSS VSS nch_mac l=30.0n w=0.14u
MM23 net37 TE VSS VSS nch_mac l=30.0n w=0.14u
MM2 net37 E VSS VSS nch_mac l=30.0n w=0.14u
MM5 qf_x clkbb net37 VSS nch_mac l=30.0n w=0.14u
MM26 qf qf_x VDD VDD pch_mac l=30.0n w=0.175u
MM25 net0245 qf VDD VDD pch_mac l=30.0n w=0.14u
MM24 qf_x clkbb net0245 VDD pch_mac l=30.0n w=0.14u
MM20 net56 net51 VDD VDD pch_mac l=30.0n w=0.17u
MM19 net11 CPN net56 VDD pch_mac l=30.0n w=0.17u
MM17 Q net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM17_2 Q net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM13 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM27 net51 qf VDD VDD pch_mac l=30.0n w=0.17u
MM12 clkb CPN VDD VDD pch_mac l=30.0n w=170.0n
MM1 qf_x clkb net88 VDD pch_mac l=30.0n w=0.14u
MM0 net88 E net92 VDD pch_mac l=30.0n w=170.0n
MM4 net92 TE VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT CKLNQD2 TE E CP Q VDD VSS
MM5 qf_x clkb net59 VSS nch_mac l=30.0n w=0.14u
MM2 net59 E VSS VSS nch_mac l=30.0n w=0.14u
MM23 net59 TE VSS VSS nch_mac l=30.0n w=0.14u
MM11 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM14 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM28 qf_x clkbb net75 VSS nch_mac l=30.0n w=0.14u
MM29 net75 qf VSS VSS nch_mac l=30.0n w=0.14u
MM30 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM9 net83 qf VSS VSS nch_mac l=30.0n w=0.14u
MM8 net39 CP net83 VSS nch_mac l=30.0n w=0.14u
MM18 Q net39 VSS VSS nch_mac l=30.0n w=0.14u 
MM18_2 Q net39 VSS VSS nch_mac l=30.0n w=0.14u 
MM4 net14 TE VDD VDD pch_mac l=30.0n w=0.17u
MM0 net18 E net14 VDD pch_mac l=30.0n w=170.0n
MM1 qf_x clkbb net18 VDD pch_mac l=30.0n w=0.14u
MM12 clkb CP VDD VDD pch_mac l=30.0n w=170.0n
MM13 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM24 qf_x clkb net30 VDD pch_mac l=30.0n w=0.14u
MM25 net30 qf VDD VDD pch_mac l=30.0n w=0.14u
MM26 qf qf_x VDD VDD pch_mac l=30.0n w=0.175u
MM7 net39 qf VDD VDD pch_mac l=30.0n w=0.185u
MM6 net39 CP VDD VDD pch_mac l=30.0n w=0.185u
MM17 Q net39 VDD VDD pch_mac l=30.0n w=0.17u 
MM17_2 Q net39 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT CKMUX2D2 I0 I1 S Z VDD VSS
MM10 Z net11 VSS VSS nch_mac l=30.0n w=0.26u 
MM10_2 Z net11 VSS VSS nch_mac l=30.0n w=0.26u 
MM7 net11 S net15 VSS nch_mac l=30.0n w=0.14u
MM6 net15 I1 VSS VSS nch_mac l=30.0n w=0.19u
MM3 net19 S VSS VSS nch_mac l=30.0n w=0.14u
MM1 net23 I0 VSS VSS nch_mac l=30.0n w=0.14u
MM5 net11 net19 net23 VSS nch_mac l=30.0n w=0.14u
MM11 Z net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM11_2 Z net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM9 net11 net19 net15 VDD pch_mac l=30.0n w=0.2u
MM8 net15 I1 VDD VDD pch_mac l=30.0n w=0.2u
MM2 net19 S VDD VDD pch_mac l=30.0n w=0.14u
MM0 net23 I0 VDD VDD pch_mac l=30.0n w=0.185u
MM4 net11 S net23 VDD pch_mac l=30.0n w=0.2u
.ENDS
.SUBCKT CKND2 I ZN VDD VSS
MM5 ZN I VSS VSS nch_mac l=30.0n w=0.25u 
MM5_2 ZN I VSS VSS nch_mac l=30.0n w=0.25u 
MM4 ZN I VDD VDD pch_mac l=30.0n w=0.32u 
MM4_2 ZN I VDD VDD pch_mac l=30.0n w=0.32u 
.ENDS
.SUBCKT CKND2D2 A1 A2 ZN VDD VSS
MM8 ZN A1 net5 VSS nch_mac l=30.0n w=0.14u 
MM8_2 ZN A1 net5 VSS nch_mac l=30.0n w=0.14u 
MM9 net5 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 net5 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 ZN A1 VDD VDD pch_mac l=30.0n w=0.165u 
MM6_2 ZN A1 VDD VDD pch_mac l=30.0n w=0.165u 
MM7 ZN A2 VDD VDD pch_mac l=30.0n w=0.165u 
MM7_2 ZN A2 VDD VDD pch_mac l=30.0n w=0.165u 
.ENDS
.SUBCKT CKXOR2D2 A1 A2 Z VDD VSS
MM9 net38 A1 net22 VSS nch_mac l=30.0n w=0.175u
MM25 net38 net18 net26 VSS nch_mac l=30.0n w=0.185u
MM7 Z net38 VSS VSS nch_mac l=30.0n w=0.18u 
MM7_2 Z net38 VSS VSS nch_mac l=30.0n w=0.18u 
MM6 net18 A1 VSS VSS nch_mac l=30.0n w=0.275u
MM1 net22 net26 VSS VSS nch_mac l=30.0n w=0.175u
MM5 net26 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM10 net38 net18 net22 VDD pch_mac l=30.0n w=0.3u
MM24 net38 A1 net26 VDD pch_mac l=30.0n w=0.3u
MM8 Z net38 VDD VDD pch_mac l=30.0n w=0.3u
MM8B Z net38 VDD VDD pch_mac l=30.0n w=0.17u
MM3 net18 A1 VDD VDD pch_mac l=30.0n w=0.12u
MM2 net22 net26 VDD VDD pch_mac l=30.0n w=245.00n
MM4 net26 A2 VDD VDD pch_mac l=30.0n w=0.3u
.ENDS
.SUBCKT DFCND2 D CP CDN Q QN VDD VSS
MM2 qf_x qf net0165 VSS nch_mac l=30.0n w=0.14u
MM3 net0165 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.25u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.25u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq net184 VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.12u
MM66 net184 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net208 VSS nch_mac l=30.0n w=140.0n
MM1 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM75 net208 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.185u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM78_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=0.295u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net0170 CDN VDD VDD pch_mac l=30.0n w=100n
MM0 mq mq_x VDD VDD pch_mac l=30.0n w=0.295u
MM61 net0170 mq VDD VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.295u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.295u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0170 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFCNQD2 D CP CDN Q VDD VSS
MM6 qf_x qf net0145 VSS nch_mac l=30.0n w=0.14u
MM7 net0145 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf clkb net0152 VSS nch_mac l=30.0n w=0.25u
MM5 net0152 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.25u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq net184 VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.12u
MM66 net184 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net208 VSS nch_mac l=30.0n w=140.0n
MM1 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM75 net208 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.185u
MM3 qf clkbb net097 VDD pch_mac l=30.0n w=0.295u
MM2 net097 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=0.295u
MM60 net0143 CDN VDD VDD pch_mac l=30.0n w=100n
MM0 mq mq_x VDD VDD pch_mac l=30.0n w=0.295u
MM61 net0143 mq VDD VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM78_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.295u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0143 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFCSND2 D CP CDN SDN Q QN VDD VSS
MM4 qf_x qf net0178 VSS nch_mac l=30.0n w=0.14u
MM5 net0178 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM2 net0176 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 net0198 mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 SDN net0176 VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.25u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.25u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq net184 VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.12u
MM66 net184 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net208 VSS nch_mac l=30.0n w=140.0n
MM49 mq SDN net0198 VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM75 net208 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.185u
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=0.295u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM3 net172 SDN VDD VDD pch_mac l=30.0n w=0.115u
MM60 net0172 CDN VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.285u
MM61 net0172 mq VDD VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM78_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.295u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.115u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0172 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT DFCSNQD2 D CP CDN SDN Q VDD VSS
MM4 qf_x qf net0178 VSS nch_mac l=30.0n w=0.14u
MM5 net0178 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM2 net0176 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 net0187 mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 SDN net0176 VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.25u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.25u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq net184 VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.12u
MM66 net184 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net208 VSS nch_mac l=30.0n w=140.0n
MM49 mq SDN net0187 VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM75 net208 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.185u
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=0.295u
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM3 net172 SDN VDD VDD pch_mac l=30.0n w=0.115u
MM60 net0161 CDN VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.285u
MM61 net0161 mq VDD VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM78_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.295u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.115u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0161 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT DFD2 D CP Q QN VDD VSS
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.27u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.27u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.175u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.18u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.175u
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=0.26u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.26u
MM60 net0132 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.26u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.175u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0132 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.175u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFKCND2 D CP CN Q QN VDD VSS
MM2 net0146 CN VSS VSS nch_mac l=30.0n w=0.135u
MM4 net172 qf_x VSS VSS nch_mac l=30.0n w=0.135u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.135u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.135u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.135u
MM66 net176 mq VSS VSS nch_mac l=30.0n w=0.135u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.135u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=0.135u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.135u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D net0146 VSS nch_mac l=30.0n w=0.135u
MM1 net090 CN VDD VDD pch_mac l=30.0n w=0.175u
MM3 net172 qf_x VDD VDD pch_mac l=30.0n w=0.185u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.175u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM60 net0143 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.185u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.185u
MM44 net090 D VDD VDD pch_mac l=30.0n w=0.175u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.185u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0143 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.185u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFKCNQD2 D CP CN Q VDD VSS
MM2 net0146 CN VSS VSS nch_mac l=30.0n w=0.25u
MM5 qf clkb net0147 VSS nch_mac l=30.0n w=0.15u
MM6 net0147 qf_x VSS VSS nch_mac l=30.0n w=0.15u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.15u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.15u
MM66 net176 mq VSS VSS nch_mac l=30.0n w=0.15u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.15u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.15u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D net0146 VSS nch_mac l=30.0n w=0.25u
MM4 qf clkbb net088 VDD pch_mac l=30.0n w=0.175u
MM1 net090 CN VDD VDD pch_mac l=30.0n w=0.175u
MM3 net088 qf_x VDD VDD pch_mac l=30.0n w=0.175u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.175u
MM60 net0128 mq VDD VDD pch_mac l=30.0n w=0.175u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net090 D VDD VDD pch_mac l=30.0n w=0.175u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0128 VDD pch_mac l=30.0n w=0.175u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.175u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFKCSND2 D CP CN SN Q QN VDD VSS
MM4 net0173 SN VSS VSS nch_mac l=30.0n w=0.14u
MM5 net212 net0173 net0146 VSS nch_mac l=30.0n w=0.12u
MM2 net0146 CN VSS VSS nch_mac l=30.0n w=0.14u
MM8 net172 qf_x VSS VSS nch_mac l=30.0n w=0.135u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.135u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.135u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.135u
MM66 net176 mq VSS VSS nch_mac l=30.0n w=0.135u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.135u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=0.135u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.135u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D net0146 VSS nch_mac l=30.0n w=0.14u
MM3 net0173 SN VDD VDD pch_mac l=30.0n w=0.12u
MM6 net0144 net0173 VDD VDD pch_mac l=30.0n w=0.215u
MM1 net090 CN VDD VDD pch_mac l=30.0n w=0.12u
MM7 net172 qf_x VDD VDD pch_mac l=30.0n w=0.185u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.215u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM60 net0163 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.185u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.185u
MM44 net090 D net0144 VDD pch_mac l=30.0n w=0.215u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.185u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0163 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.185u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFKSND2 D CP SN Q QN VDD VSS
MM4 net0173 SN VSS VSS nch_mac l=30.0n w=0.14u
MM5 net212 net0173 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net172 qf_x VSS VSS nch_mac l=30.0n w=0.135u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.135u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.135u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.135u
MM66 net176 mq VSS VSS nch_mac l=30.0n w=0.135u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.135u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=0.135u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.135u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.14u
MM3 net0173 SN VDD VDD pch_mac l=30.0n w=0.12u
MM6 net0144 net0173 VDD VDD pch_mac l=30.0n w=170.0n
MM7 net172 qf_x VDD VDD pch_mac l=30.0n w=0.185u
MM45 mq_x clkbb net212 VDD pch_mac l=30.0n w=0.215u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM60 net0153 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.185u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.185u
MM44 net212 D net0144 VDD pch_mac l=30.0n w=0.17u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.185u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0153 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.185u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFMD2 DA DB SA CP Q QN VDD VSS
MM8 net0184 DA VSS VSS nch_mac l=30.0n w=0.17u
MM4 net0176 SA VSS VSS nch_mac l=30.0n w=0.14u
MM9 net212 SA net0184 VSS nch_mac l=30.0n w=170.0n
MM2 net0231 DB VSS VSS nch_mac l=30.0n w=0.17u
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.27u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.27u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.175u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 net0176 net0231 VSS nch_mac l=30.0n w=0.17u
MM7 net0119 DA VDD VDD pch_mac l=30.0n w=0.27u
MM3 net0176 SA VDD VDD pch_mac l=30.0n w=0.27u
MM6 net0231 DB VDD VDD pch_mac l=30.0n w=0.27u
MM1 net090 net0176 net0119 VDD pch_mac l=30.0n w=0.27u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.24u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.26u
MM60 net0171 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.175u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net090 SA net0231 VDD pch_mac l=30.0n w=0.27u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.25u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0171 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.175u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=135.0n
.ENDS
.SUBCKT DFMQD2 DA DB SA CP Q VDD VSS
MM8 net0184 DA VSS VSS nch_mac l=30.0n w=0.17u
MM12 qf clkb net0177 VSS nch_mac l=30.0n w=0.14u
MM4 net0176 SA VSS VSS nch_mac l=30.0n w=0.14u
MM13 net0177 qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM9 net212 SA net0184 VSS nch_mac l=30.0n w=170.0n
MM2 net0146 DB VSS VSS nch_mac l=30.0n w=0.17u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.14u
MM66 net176 mq VSS VSS nch_mac l=30.0n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.25u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.175u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 net0176 net0146 VSS nch_mac l=30.0n w=0.17u
MM7 net0119 DA VDD VDD pch_mac l=30.0n w=0.27u
MM3 net0176 SA VDD VDD pch_mac l=30.0n w=0.27u
MM6 net0146 DB VDD VDD pch_mac l=30.0n w=0.27u
MM1 net090 net0176 net0119 VDD pch_mac l=30.0n w=0.27u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.24u
MM60 net0171 mq VDD VDD pch_mac l=30.0n w=0.18u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.18u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.3u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net090 SA net0146 VDD pch_mac l=30.0n w=0.27u
MM10 net0116 qf_x VDD VDD pch_mac l=30.0n w=0.18u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0171 VDD pch_mac l=30.0n w=0.18u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.18u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=135.0n
MM11 qf clkbb net0116 VDD pch_mac l=30.0n w=0.18u
.ENDS
.SUBCKT DFNCND2 D CPN CDN Q QN VDD VSS
MM2 qf_x qf net0165 VSS nch_mac l=30.0n w=0.14u
MM3 net0165 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.25u
MM67 net172 clkbb qf VSS nch_mac l=30.0n w=0.25u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq net184 VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkb net176 VSS nch_mac l=30.0n w=0.12u
MM66 net184 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkbb net212 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net208 VSS nch_mac l=30.0n w=140.0n
MM1 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=0.14u
MM75 net208 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.185u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM78_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkb net103 VDD pch_mac l=30.0n w=0.295u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net0170 CDN VDD VDD pch_mac l=30.0n w=100n
MM0 mq mq_x VDD VDD pch_mac l=30.0n w=0.295u
MM61 net0170 mq VDD VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.295u
MM68 net172 clkb qf VDD pch_mac l=30.0n w=0.295u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkbb net0170 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFNCSND2 D CPN CDN SDN Q QN VDD VSS
MM4 qf_x qf net0178 VSS nch_mac l=30.0n w=0.14u
MM5 net0178 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM2 net0176 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 net0198 mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 SDN net0176 VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.25u
MM67 net172 clkbb qf VSS nch_mac l=30.0n w=0.25u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq net184 VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkb net176 VSS nch_mac l=30.0n w=0.12u
MM66 net184 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkbb net212 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net208 VSS nch_mac l=30.0n w=140.0n
MM49 mq SDN net0198 VSS nch_mac l=30.0n w=0.14u
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=0.14u
MM75 net208 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.185u
MM45 mq_x clkb net103 VDD pch_mac l=30.0n w=0.295u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM3 net172 SDN VDD VDD pch_mac l=30.0n w=0.115u
MM60 net0172 CDN VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.285u
MM61 net0172 mq VDD VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM78_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.295u
MM68 net172 clkb qf VDD pch_mac l=30.0n w=0.115u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkbb net0172 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT DFND2 D CPN Q QN VDD VSS
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.27u
MM67 net172 clkbb qf VSS nch_mac l=30.0n w=0.27u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkbb net212 VSS nch_mac l=30.0n w=0.175u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.18u
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.175u
MM45 mq_x clkb net103 VDD pch_mac l=30.0n w=0.26u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.26u
MM60 net0132 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.26u
MM68 net172 clkb qf VDD pch_mac l=30.0n w=0.175u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkbb net0132 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.175u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFNSND2 D CPN SDN Q QN VDD VSS
MM2 net0176 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 net0162 mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 SDN net0176 VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.22u
MM67 net172 clkbb qf VSS nch_mac l=30.0n w=0.22u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq VSS VSS nch_mac l=30.0n w=0.14u
MM64 mq_x clkb net176 VSS nch_mac l=30.0n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkbb net212 VSS nch_mac l=30.0n w=0.14u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq SDN net0162 VSS nch_mac l=30.0n w=0.14u
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=140.0n
MM45 mq_x clkb net103 VDD pch_mac l=30.0n w=200n
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM3 net172 SDN VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.31u
MM61 net0144 mq VDD VDD pch_mac l=30.0n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.2u
MM68 net172 clkb qf VDD pch_mac l=30.0n w=0.11u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkbb net0144 VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.31u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.2u
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT DFQD2 D CP Q VDD VSS
MM2 qf clkb net0136 VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.175u
MM3 net0136 qf_x VSS VSS nch_mac l=30.0n w=0.175u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.175u
MM66 net176 mq VSS VSS nch_mac l=30.0n w=0.175u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.175u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.175u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=0.175u
MM0 net086 qf_x VDD VDD pch_mac l=30.0n w=0.175u
MM1 qf clkbb net086 VDD pch_mac l=30.0n w=0.175u
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=0.26u
MM60 net0118 mq VDD VDD pch_mac l=30.0n w=0.175u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.26u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0118 VDD pch_mac l=30.0n w=0.175u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.175u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT DFSND2 D CP SDN Q QN VDD VSS
MM2 net0176 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 net0162 mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 SDN net0176 VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.22u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.22u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq VSS VSS nch_mac l=30.0n w=0.14u
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.195u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.195u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq SDN net0162 VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=140.0n
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=200n
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM3 net172 SDN VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.31u
MM61 net0144 mq VDD VDD pch_mac l=30.0n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.2u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.11u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0144 VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.31u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.2u
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT DFSNQD2 D CP SDN Q VDD VSS
MM2 net0176 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 net0162 mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM73 net172 SDN net0176 VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.22u
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.22u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net176 mq VSS VSS nch_mac l=30.0n w=0.14u
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=0.195u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.195u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq SDN net0162 VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.14u
MM47 net212 D VSS VSS nch_mac l=30.0n w=140.0n
MM45 mq_x clkbb net103 VDD pch_mac l=30.0n w=200n
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM3 net172 SDN VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.31u
MM61 net0144 mq VDD VDD pch_mac l=30.0n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net103 D VDD VDD pch_mac l=30.0n w=0.2u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.11u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0144 VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.31u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.2u
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT EDFCND2 D E CP CDN Q QN VDD VSS
MM14 net0215 CDN VSS VSS nch_mac l=30.0n w=0.195u
MM15 qf_x qf net0215 VSS nch_mac l=30.0n w=0.14u
MM11 net0209 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM13 net0201 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM8 net0184 D VSS VSS nch_mac l=30.0n w=0.175u
MM4 net0176 E VSS VSS nch_mac l=30.0n w=0.22u
MM9 net212 E net0184 VSS nch_mac l=30.0n w=0.175u
MM2 net0146 net172 VSS VSS nch_mac l=30.0n w=0.175u
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.195u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=275.00n
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.195u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq net0201 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.17u
MM76 qf_x qf net0209 VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.27u
MM47 net212 net0176 net0146 VSS nch_mac l=30.0n w=0.175u
MM0 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u
MM0B qf_x CDN VDD VDD pch_mac l=30.0n w=0.26u
MM12 net0199 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM7 net0184 D VDD VDD pch_mac l=30.0n w=0.27u
MM3 net0176 E VDD VDD pch_mac l=30.0n w=0.12u
MM6 net0144 net172 VDD VDD pch_mac l=30.0n w=0.27u
MM1 net090 net0176 net0184 VDD pch_mac l=30.0n w=0.27u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.265u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.26u
MM60 net0199 mq VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.275u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM44 net090 E net0144 VDD pch_mac l=30.0n w=0.27u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0199 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=135.0n
.ENDS
.SUBCKT EDFCNQD2 D E CP CDN Q VDD VSS
MM15 qf_x qf net0204 VSS nch_mac l=30.0n w=0.14u
MM11 net0196 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM14 net0204 CDN VSS VSS nch_mac l=30.0n w=0.195u
MM13 net0201 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM8 net0184 D VSS VSS nch_mac l=30.0n w=0.175u
MM4 net0176 E VSS VSS nch_mac l=30.0n w=0.22u
MM9 net212 E net0184 VSS nch_mac l=30.0n w=0.175u
MM2 net0146 net172 VSS VSS nch_mac l=30.0n w=0.175u
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.195u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=275.00n
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.195u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq net0201 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.17u
MM76 qf_x qf net0196 VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.27u
MM47 net212 net0176 net0146 VSS nch_mac l=30.0n w=0.175u
MM0 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u
MM0B qf_x CDN VDD VDD pch_mac l=30.0n w=0.26u
MM12 net0199 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM7 net0184 D VDD VDD pch_mac l=30.0n w=0.27u
MM3 net0176 E VDD VDD pch_mac l=30.0n w=0.12u
MM6 net0144 net172 VDD VDD pch_mac l=30.0n w=0.27u
MM1 net090 net0176 net0184 VDD pch_mac l=30.0n w=0.27u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.265u
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.26u
MM60 net0199 mq VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.275u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM44 net090 E net0144 VDD pch_mac l=30.0n w=0.27u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0199 VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=135.0n
.ENDS
.SUBCKT EDFD2 D E CP Q QN VDD VSS
MM8 net0184 D VSS VSS nch_mac l=30.0n w=0.175u
MM4 net0176 E VSS VSS nch_mac l=30.0n w=0.25u
MM9 net212 E net0184 VSS nch_mac l=30.0n w=0.175u
MM2 net0146 net172 VSS VSS nch_mac l=30.0n w=0.175u
MM16 net172 qf_x VSS VSS nch_mac l=30.0n w=0.275u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=275.00n
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.275u
MM69 QN net172 VSS VSS nch_mac l=30.0n w=0.275u 
MM69_2 QN net172 VSS VSS nch_mac l=30.0n w=0.275u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.17u
MM14 qf_x qf VSS VSS nch_mac l=30.0n w=0.14u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.27u
MM47 net212 net0176 net0146 VSS nch_mac l=30.0n w=0.175u
MM7 net0184 D VDD VDD pch_mac l=30.0n w=0.27u
MM3 net0176 E VDD VDD pch_mac l=30.0n w=0.12u
MM6 net0144 net172 VDD VDD pch_mac l=30.0n w=0.27u
MM1 net090 net0176 net0184 VDD pch_mac l=30.0n w=0.27u
MM15 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.265u
MM70 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net172 VDD VDD pch_mac l=30.0n w=0.17u 
MM60 net0173 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.275u
MM13 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u
MM44 net090 E net0144 VDD pch_mac l=30.0n w=0.27u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0173 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=135.0n
.ENDS
.SUBCKT EDFQD2 D E CP Q VDD VSS
MM8 net0184 D VSS VSS nch_mac l=30.0n w=0.175u
MM4 net0176 E VSS VSS nch_mac l=30.0n w=0.25u
MM9 net212 E net0184 VSS nch_mac l=30.0n w=0.175u
MM2 net0146 net172 VSS VSS nch_mac l=30.0n w=0.175u
MM73 net172 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=275.00n
MM67 net172 clkb qf VSS nch_mac l=30.0n w=0.275u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM64 mq_x clkbb net176 VSS nch_mac l=30.0n w=100n
MM66 net176 mq VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net212 VSS nch_mac l=30.0n w=0.17u
MM14 qf_x qf VSS VSS nch_mac l=30.0n w=0.14u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.27u
MM47 net212 net0176 net0146 VSS nch_mac l=30.0n w=0.175u
MM7 net0184 D VDD VDD pch_mac l=30.0n w=0.27u
MM3 net0176 E VDD VDD pch_mac l=30.0n w=0.12u
MM6 net0144 net172 VDD VDD pch_mac l=30.0n w=0.27u
MM1 net090 net0176 net0184 VDD pch_mac l=30.0n w=0.27u
MM45 mq_x clkbb net090 VDD pch_mac l=30.0n w=0.265u
MM74 net172 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net0173 mq VDD VDD pch_mac l=30.0n w=100n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.275u
MM13 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u
MM44 net090 E net0144 VDD pch_mac l=30.0n w=0.27u
MM68 net172 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net0173 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=135.0n
.ENDS
.SUBCKT FA1D2 A B CI S CO VDD VSS
MM22 net172 net148 net184 VSS nch_mac l=30n w=0.14u
MM21 net184 B VSS VSS nch_mac l=30n w=0.14u
MM34 net184 CI VSS VSS nch_mac l=30n w=0.14u
MM38 net176 CI VSS VSS nch_mac l=30n w=0.14u
MM15 net172 A net144 VSS nch_mac l=30n w=0.14u
MM14 S net172 VSS VSS nch_mac l=30n w=0.14u 
MM14_2 S net172 VSS VSS nch_mac l=30n w=0.14u 
MM13 net160 A VSS VSS nch_mac l=30n w=0.275u
MM12 net160 B VSS VSS nch_mac l=30n w=0.275u
MM11 net148 CI net160 VSS nch_mac l=30n w=140n
MM6 CO net148 VSS VSS nch_mac l=30n w=0.14u 
MM6_2 CO net148 VSS VSS nch_mac l=30n w=0.14u 
MM4 net148 A net140 VSS nch_mac l=30n w=0.275u
MM37 net144 B net176 VSS nch_mac l=30n w=140n
MM5 net140 B VSS VSS nch_mac l=30n w=0.275u
MM33 net184 A VSS VSS nch_mac l=30n w=0.14u
MM31 net239 CI VDD VDD pch_mac l=30n w=0.17u
MM32 net172 net148 net239 VDD pch_mac l=30n w=0.17u
MM25 net239 B VDD VDD pch_mac l=30n w=0.17u
MM35 net226 B net238 VDD pch_mac l=30n w=0.17u
MM30 net239 A VDD VDD pch_mac l=30n w=0.17u
MM17 S net172 VDD VDD pch_mac l=30n w=0.17u 
MM17_2 S net172 VDD VDD pch_mac l=30n w=0.17u 
MM36 net172 A net226 VDD pch_mac l=30n w=170n
MM10 net148 CI net211 VDD pch_mac l=30n w=0.21u
MM28 net238 CI VDD VDD pch_mac l=30n w=0.17u
MM8 net211 B VDD VDD pch_mac l=30n w=0.17u
MM9 net211 A VDD VDD pch_mac l=30n w=0.17u
MM2 net198 B VDD VDD pch_mac l=30n w=0.21u
MM7 CO net148 VDD VDD pch_mac l=30n w=0.17u 
MM7_2 CO net148 VDD VDD pch_mac l=30n w=0.17u 
MM3 net148 A net198 VDD pch_mac l=30n w=0.21u
.ENDS
.SUBCKT FA1OPTCD2 A B CI S CO VDD VSS
MM22 net172 net148 net184 VSS nch_mac l=30n w=0.14u
MM21 net184 B VSS VSS nch_mac l=30n w=0.14u
MM34 net184 CI VSS VSS nch_mac l=30n w=0.14u
MM38 net176 CI VSS VSS nch_mac l=30n w=0.14u
MM15 net172 A net144 VSS nch_mac l=30n w=0.14u
MM14 S net172 VSS VSS nch_mac l=30n w=0.14u 
MM14_2 S net172 VSS VSS nch_mac l=30n w=0.14u 
MM13 net160 A VSS VSS nch_mac l=30n w=0.14u 
MM13_2 net160 A VSS VSS nch_mac l=30n w=0.14u 
MM13_3 net160 A VSS VSS nch_mac l=30n w=0.14u 
MM12 net160 B VSS VSS nch_mac l=30n w=0.14u 
MM12_2 net160 B VSS VSS nch_mac l=30n w=0.14u 
MM12_3 net160 B VSS VSS nch_mac l=30n w=0.14u 
MM11 net148 CI net160 VSS nch_mac l=30n w=0.14u 
MM11_2 net148 CI net160 VSS nch_mac l=30n w=0.14u 
MM6 CO net148 VSS VSS nch_mac l=30n w=0.14u 
MM6_2 CO net148 VSS VSS nch_mac l=30n w=0.14u 
MM4 net148 A net140 VSS nch_mac l=30n w=0.14u
MM37 net144 B net176 VSS nch_mac l=30n w=140n
MM5 net140 B VSS VSS nch_mac l=30n w=0.14u
MM33 net184 A VSS VSS nch_mac l=30n w=0.14u
MM31 net239 CI VDD VDD pch_mac l=30n w=0.17u
MM32 net172 net148 net239 VDD pch_mac l=30n w=0.17u
MM25 net239 B VDD VDD pch_mac l=30n w=0.17u
MM35 net226 B net238 VDD pch_mac l=30n w=0.17u
MM30 net239 A VDD VDD pch_mac l=30n w=0.17u
MM17 S net172 VDD VDD pch_mac l=30n w=0.17u 
MM17_2 S net172 VDD VDD pch_mac l=30n w=0.17u 
MM36 net172 A net226 VDD pch_mac l=30n w=170n
MM10 net148 CI net211 VDD pch_mac l=30n w=0.17u 
MM10_2 net148 CI net211 VDD pch_mac l=30n w=0.17u 
MM28 net238 CI VDD VDD pch_mac l=30n w=0.17u
MM8 net211 B VDD VDD pch_mac l=30n w=0.17u 
MM8_2 net211 B VDD VDD pch_mac l=30n w=0.17u 
MM8_3 net211 B VDD VDD pch_mac l=30n w=0.17u 
MM9 net211 A VDD VDD pch_mac l=30n w=0.17u 
MM9_2 net211 A VDD VDD pch_mac l=30n w=0.17u 
MM9_3 net211 A VDD VDD pch_mac l=30n w=0.17u 
MM2 net198 B VDD VDD pch_mac l=30n w=0.17u
MM7 CO net148 VDD VDD pch_mac l=30n w=0.17u 
MM7_2 CO net148 VDD VDD pch_mac l=30n w=0.17u 
MM3 net148 A net198 VDD pch_mac l=30n w=0.17u
.ENDS
.SUBCKT FA1OPTSD2 A B CI S CO VDD VSS
MM9 net111 A VDD VDD pch_mac l=30n w=0.17u 
MM9_2 net111 A VDD VDD pch_mac l=30n w=0.17u 
MM36 net160 A net130 VDD pch_mac l=30n w=170n
MM10 net172 CI net111 VDD pch_mac l=30n w=0.17u 
MM10_2 net172 CI net111 VDD pch_mac l=30n w=0.17u 
MM30 net115 A VDD VDD pch_mac l=30n w=0.17u 
MM30_2 net115 A VDD VDD pch_mac l=30n w=0.17u 
MM30_3 net115 A VDD VDD pch_mac l=30n w=0.17u 
MM25 net115 B VDD VDD pch_mac l=30n w=0.17u 
MM25_2 net115 B VDD VDD pch_mac l=30n w=0.17u 
MM25_3 net115 B VDD VDD pch_mac l=30n w=0.17u 
MM8 net111 B VDD VDD pch_mac l=30n w=0.17u 
MM8_2 net111 B VDD VDD pch_mac l=30n w=0.17u 
MM32 net160 net172 net115 VDD pch_mac l=30n w=0.17u 
MM32_2 net160 net172 net115 VDD pch_mac l=30n w=0.17u 
MM35 net130 B net106 VDD pch_mac l=30n w=0.17u
MM7 CO net172 VDD VDD pch_mac l=30n w=0.17u 
MM7_2 CO net172 VDD VDD pch_mac l=30n w=0.17u 
MM3 net172 A net154 VDD pch_mac l=30n w=0.17u
MM2 net154 B VDD VDD pch_mac l=30n w=0.17u
MM28 net106 CI VDD VDD pch_mac l=30n w=0.17u
MM31 net115 CI VDD VDD pch_mac l=30n w=0.17u 
MM31_2 net115 CI VDD VDD pch_mac l=30n w=0.17u 
MM31_3 net115 CI VDD VDD pch_mac l=30n w=0.17u 
MM17 S net160 VDD VDD pch_mac l=30n w=0.17u 
MM17_2 S net160 VDD VDD pch_mac l=30n w=0.17u 
MM34 net188 CI VSS VSS nch_mac l=30n w=0.14u 
MM34_2 net188 CI VSS VSS nch_mac l=30n w=0.14u 
MM34_3 net188 CI VSS VSS nch_mac l=30n w=0.14u 
MM12 net192 B VSS VSS nch_mac l=30n w=0.14u 
MM12_2 net192 B VSS VSS nch_mac l=30n w=0.14u 
MM13 net192 A VSS VSS nch_mac l=30n w=0.14u 
MM13_2 net192 A VSS VSS nch_mac l=30n w=0.14u 
MM38 net204 CI VSS VSS nch_mac l=30n w=0.14u
MM6 CO net172 VSS VSS nch_mac l=30n w=0.14u 
MM6_2 CO net172 VSS VSS nch_mac l=30n w=0.14u 
MM33 net188 A VSS VSS nch_mac l=30n w=0.14u 
MM33_2 net188 A VSS VSS nch_mac l=30n w=0.14u 
MM33_3 net188 A VSS VSS nch_mac l=30n w=0.14u 
MM4 net172 A net164 VSS nch_mac l=30n w=0.14u
MM22 net160 net172 net188 VSS nch_mac l=30n w=0.14u 
MM22_2 net160 net172 net188 VSS nch_mac l=30n w=0.14u 
MM37 net168 B net204 VSS nch_mac l=30n w=140n
MM5 net164 B VSS VSS nch_mac l=30n w=0.14u
MM15 net160 A net168 VSS nch_mac l=30n w=0.14u
MM14 S net160 VSS VSS nch_mac l=30n w=0.14u 
MM14_2 S net160 VSS VSS nch_mac l=30n w=0.14u 
MM21 net188 B VSS VSS nch_mac l=30n w=0.14u 
MM21_2 net188 B VSS VSS nch_mac l=30n w=0.14u 
MM21_3 net188 B VSS VSS nch_mac l=30n w=0.14u 
MM11 net172 CI net192 VSS nch_mac l=30n w=0.14u 
MM11_2 net172 CI net192 VSS nch_mac l=30n w=0.14u 
.ENDS
.SUBCKT GAN2D2 A1 A2 Z VDD VSS
MM9 net14 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net26 A1 net14 VSS nch_mac l=30.0n w=0.14u
MM5 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net26 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM7 net26 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM4 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT GAOI21D2 A1 A2 B ZN VDD VSS
MM5 ZN A1 net027 VSS nch_mac l=30.0n w=0.14u
MM4 net027 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM2 net7 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM1 ZN A1 net7 VSS nch_mac l=30.0n w=0.14u
MM0 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net30 B VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 net30 B VDD VDD pch_mac l=30.0n w=0.17u 
MM6 ZN A2 net30 VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN A2 net30 VDD pch_mac l=30.0n w=0.17u 
MM3 ZN A1 net30 VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN A1 net30 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT GBUFFD2 I Z VDD VSS
MM26 VSS I VSS VSS nch_mac l=30.0n w=0.14u
MM0 Z net9 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net9 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net9 I VSS VSS nch_mac l=30.0n w=0.14u
MM24 VDD I VDD VDD pch_mac l=30.0n w=170.0n
MM1 Z net9 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net9 VDD VDD pch_mac l=30.0n w=0.17u 
MM4 net9 I VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GINVD2 I ZN VDD VSS
MM1 ZN I VSS VSS nch_mac l=30.0n w=0.14u 
MM1_2 ZN I VSS VSS nch_mac l=30.0n w=0.14u 
MM0 ZN I VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 ZN I VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT GMUX2D2 I0 I1 S Z VDD VSS
MM6 net57 I1 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 net57 I1 VSS VSS nch_mac l=30.0n w=0.14u 
MM9 net85 S VSS VSS nch_mac l=30.0n w=0.14u
MM2 net62 I0 VSS VSS nch_mac l=30.0n w=0.14u
MM7 net53 S net57 VSS nch_mac l=30.0n w=0.14u
MM12 Z net53 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Z net53 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net53 net85 net62 VSS nch_mac l=30.0n w=0.14u
MM14 net93 I1 VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 net93 I1 VDD VDD pch_mac l=30.0n w=0.17u 
MM8 net85 S VDD VDD pch_mac l=30.0n w=0.17u
MM13 Z net53 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Z net53 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 net53 S net97 VDD pch_mac l=30.0n w=0.17u
MM3 net97 I0 VDD VDD pch_mac l=30.0n w=0.17u
MM5 net53 net85 net93 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GMUX2ND2 I0 I1 S ZN VDD VSS
MM15 ZN net103 VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 ZN net103 VSS VSS nch_mac l=30.0n w=0.14u 
MM11 net103 net87 VSS VSS nch_mac l=30.0n w=140.0n
MM0 net87 net83 net63 VSS nch_mac l=30.0n w=0.14u
MM2 net63 I0 VSS VSS nch_mac l=30.0n w=0.14u
MM7 net87 S net59 VSS nch_mac l=30.0n w=0.14u
MM6 net59 I1 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net83 S VSS VSS nch_mac l=30.0n w=0.14u
MM14 ZN net103 VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 ZN net103 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 net103 net87 VDD VDD pch_mac l=30.0n w=0.17u
MM1 net87 S net95 VDD pch_mac l=30.0n w=0.17u
MM8 net83 S VDD VDD pch_mac l=30.0n w=0.17u
MM3 net95 I0 VDD VDD pch_mac l=30.0n w=0.17u
MM4 net84 I1 VDD VDD pch_mac l=30.0n w=0.17u
MM5 net87 net83 net84 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GND2D2 A1 A2 ZN VDD VSS
MM0 net33 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM3 ZN A1 net33 VSS nch_mac l=30.0n w=0.14u
MM7 net28 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM6 ZN A1 net28 VSS nch_mac l=30.0n w=0.14u
MM2 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT GND3D2 A1 A2 A3 ZN VDD VSS
MM7 net33 A2 net61 VSS nch_mac l=30.0n w=0.14u
MM8 ZN A1 net33 VSS nch_mac l=30.0n w=0.14u
MM2 net41 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM1 net46 A2 net41 VSS nch_mac l=30.0n w=0.14u
MM0 ZN A1 net46 VSS nch_mac l=30.0n w=0.14u
MM6 net61 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM4 ZN A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM5 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM5_2 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT GNR2D2 A1 A2 ZN VDD VSS
MM1 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM1_2 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM3 ZN A2 net45 VDD pch_mac l=30.0n w=0.17u
MM6 net37 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM4 ZN A2 net37 VDD pch_mac l=30.0n w=0.17u
MM2 net45 A1 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GNR3D2 A1 A2 A3 ZN VDD VSS
MM0 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM3 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM1 ZN A3 VSS VSS nch_mac l=30.0n w=0.14u 
MM1_2 ZN A3 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net56 A2 net44 VDD pch_mac l=30.0n w=0.17u 
MM6_2 net56 A2 net44 VDD pch_mac l=30.0n w=0.17u 
MM4 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN A1 net56 VDD pch_mac l=30.0n w=0.17u 
MM2 net44 A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 net44 A3 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT GOAI21D2 A1 A2 B ZN VDD VSS
MM3 net30 B VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 net30 B VSS VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A2 net30 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A2 net30 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A1 net30 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A1 net30 VSS nch_mac l=30.0n w=0.14u 
MM4 ZN A1 net031 VDD pch_mac l=30.0n w=0.17u
MM5 net031 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM59 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM59_2 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM0 ZN A1 net14 VDD pch_mac l=30.0n w=170.0n
MM1 net14 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GOR2D2 A1 A2 Z VDD VSS
MM0 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM8 net26 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net26 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM1 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net26 A1 net13 VDD pch_mac l=30.0n w=0.17u
MM7 net13 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GXNR2D2 A1 A2 ZN VDD VSS
MM3 net37 net62 net49 VSS nch_mac l=30.0n w=0.14u
MM1 net49 net40 VSS VSS nch_mac l=30.0n w=0.14u
MM6 ZN net37 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 ZN net37 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net40 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 net40 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM17 net40 A1 net37 VSS nch_mac l=30.0n w=0.14u
MM8 net62 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM15 net37 A1 net80 VDD pch_mac l=30.0n w=0.17u
MM14 net80 net40 VDD VDD pch_mac l=30.0n w=170.0n
MM7 ZN net37 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 ZN net37 VDD VDD pch_mac l=30.0n w=0.17u 
MM2 net40 A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 net40 A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net40 net62 net37 VDD pch_mac l=30.0n w=0.17u
MM9 net62 A1 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT GXOR2D2 A1 A2 Z VDD VSS
MM1 net56 net57 VSS VSS nch_mac l=30.0n w=0.14u
MM3 net60 A1 net56 VSS nch_mac l=30.0n w=0.14u
MM8 net34 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM0 net57 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 net57 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 Z net60 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 Z net60 VSS VSS nch_mac l=30.0n w=0.14u 
MM17 net60 net34 net57 VSS nch_mac l=30.0n w=0.14u
MM15 net60 net34 net77 VDD pch_mac l=30.0n w=0.17u
MM14 net77 net57 VDD VDD pch_mac l=30.0n w=170.0n
MM7 Z net60 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 Z net60 VDD VDD pch_mac l=30.0n w=0.17u 
MM9 net34 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM2 net57 A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 net57 A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net60 A1 net57 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT HA1D2 A B S CO VDD VSS
MM18 net92 A VDD VDD pch_mac l=30.0n w=0.17u
MM18B net92 A VDD VDD pch_mac l=30.0n w=0.17u
MM17 net104 B VDD VDD pch_mac l=30.0n w=0.17u
MM16 net104 A VDD VDD pch_mac l=30.0n w=0.17u
MM13 CO net104 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 CO net104 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net88 net92 VDD VDD pch_mac l=30.0n w=0.17u
MM4 net88 net124 net129 VDD pch_mac l=30.0n w=0.26u
MM7 net92 B net129 VDD pch_mac l=30.0n w=0.26u
MM9 S net129 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_2 S net129 VDD VDD pch_mac l=30.0n w=0.17u 
MM11 net124 B VDD VDD pch_mac l=30.0n w=0.17u
MM1 net92 A VSS VSS nch_mac l=30.0n w=0.26u 
MM1_2 net92 A VSS VSS nch_mac l=30.0n w=0.26u 
MM2 net88 net92 VSS VSS nch_mac l=30.0n w=0.26u
MM5 net88 B net129 VSS nch_mac l=30.0n w=0.26u
MM6 net92 net124 net129 VSS nch_mac l=30.0n w=0.26u
MM8 S net129 VSS VSS nch_mac l=30.0n w=0.14u 
MM8_2 S net129 VSS VSS nch_mac l=30.0n w=0.14u 
MM10 net124 B VSS VSS nch_mac l=30.0n w=0.14u
MM12 CO net104 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 CO net104 VSS VSS nch_mac l=30.0n w=0.14u 
MM14 net104 A net113 VSS nch_mac l=30.0n w=0.27u
MM15 net113 B VSS VSS nch_mac l=30.0n w=0.27u
.ENDS
.SUBCKT IAO21D2 A1 A2 B ZN VDD VSS
MM6 ZN net27 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 ZN net27 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 ZN B VSS VSS nch_mac l=30.0n w=0.14u 
MM3 net27 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM4 net27 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM2 net045 net27 VDD VDD pch_mac l=30.0n w=0.17u
MM1 net27 A1 net43 VDD pch_mac l=30.0n w=0.17u
MM0 net43 A2 VDD VDD pch_mac l=30.0n w=170.0n
MM7 net39 net27 VDD VDD pch_mac l=30.0n w=0.17u
MM8 ZN B net39 VDD pch_mac l=30.0n w=0.17u
MM9 ZN B net045 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT IAO22D2 A1 A2 B1 B2 ZN VDD VSS
MM13 net52 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM13_2 net52 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM12 ZN net36 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 ZN net36 VSS VSS nch_mac l=30.0n w=0.14u 
MM9 ZN B1 net52 VSS nch_mac l=30.0n w=0.14u 
MM9_2 ZN B1 net52 VSS nch_mac l=30.0n w=0.14u 
MM15 net36 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM18 net36 A1 VSS VSS nch_mac l=30.0n w=140n
MM10 net64 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM10_2 net64 B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM11 ZN net36 net64 VDD pch_mac l=30.0n w=0.17u 
MM11_2 ZN net36 net64 VDD pch_mac l=30.0n w=0.17u 
MM2 net64 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 net64 B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net59 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM17 net36 A1 net59 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT IND2D2 A1 B1 ZN VDD VSS
MM7 net024 B1 VSS VSS nch_mac l=30.0n w=0.14u
MM6 ZN net052 net024 VSS nch_mac l=30.0n w=0.14u
MM4 ZN net052 net036 VSS nch_mac l=30.0n w=0.14u
MM5 net036 B1 VSS VSS nch_mac l=30.0n w=0.14u
MM1 net052 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM2 ZN B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 ZN B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 ZN net052 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN net052 VDD VDD pch_mac l=30.0n w=0.17u 
MM0 net052 A1 VDD VDD pch_mac l=30.0n w=170.0n
.ENDS
.SUBCKT IND3D2 A1 B1 B2 ZN VDD VSS
MM1 net37 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM4 ZN B2 net57 VSS nch_mac l=30.0n w=0.14u 
MM4_2 ZN B2 net57 VSS nch_mac l=30.0n w=0.14u 
MM5 net57 B1 net53 VSS nch_mac l=30.0n w=0.14u 
MM5_2 net57 B1 net53 VSS nch_mac l=30.0n w=0.14u 
MM7 net53 net37 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net53 net37 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net37 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM2 ZN B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 ZN B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 ZN B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 ZN net37 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN net37 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT IND4D2 A1 B1 B2 B3 ZN VDD VSS
MM0 net50 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM8 ZN net50 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_2 ZN net50 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 ZN B3 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN B3 VDD VDD pch_mac l=30.0n w=0.17u 
MM2 ZN B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 ZN B2 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 ZN B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 ZN B1 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 net50 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net64 net50 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 net64 net50 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net60 B1 net64 VSS nch_mac l=30.0n w=0.14u 
MM7_2 net60 B1 net64 VSS nch_mac l=30.0n w=0.14u 
MM5 net59 B2 net60 VSS nch_mac l=30.0n w=0.14u 
MM5_2 net59 B2 net60 VSS nch_mac l=30.0n w=0.14u 
MM4 ZN B3 net59 VSS nch_mac l=30.0n w=0.14u 
MM4_2 ZN B3 net59 VSS nch_mac l=30.0n w=0.14u 
.ENDS
.SUBCKT INR2D2 A1 B1 ZN VDD VSS
MM1 net37 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM2 ZN B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM3 ZN net37 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 ZN net37 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net034 net37 VDD VDD pch_mac l=30.0n w=170.0n
MM0 net37 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM7 ZN B1 net034 VDD pch_mac l=30.0n w=0.17u
MM4 ZN B1 net29 VDD pch_mac l=30.0n w=0.17u
MM5 net29 net37 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT INR3D2 A1 B1 B2 ZN VDD VSS
MM1 net74 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM7 ZN B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 ZN B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 ZN B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM3 ZN net74 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 ZN net74 VSS VSS nch_mac l=30.0n w=0.14u 
MM10 ZN B2 net54 VDD pch_mac l=30.0n w=0.17u
MM9 net54 B1 net50 VDD pch_mac l=30.0n w=0.17u
MM8 net50 net74 VDD VDD pch_mac l=30.0n w=0.17u
MM0 net74 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM6 net37 net74 VDD VDD pch_mac l=30.0n w=170.0n
MM4 ZN B2 net34 VDD pch_mac l=30.0n w=0.17u
MM5 net34 B1 net37 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT INR4D2 A1 B1 B2 B3 ZN VDD VSS
MM9 ZN B3 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 ZN B3 VSS VSS nch_mac l=30.0n w=0.14u 
MM1 net50 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM3 ZN net50 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 ZN net50 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 ZN B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 ZN B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 ZN B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net50 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM8 net69 net50 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_2 net69 net50 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_3 net69 net50 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_4 net69 net50 VDD VDD pch_mac l=30.0n w=0.17u 
MM5 net65 B2 net66 VDD pch_mac l=30.0n w=0.17u 
MM5_2 net65 B2 net66 VDD pch_mac l=30.0n w=0.17u 
MM5_3 net65 B2 net66 VDD pch_mac l=30.0n w=0.17u 
MM5_4 net65 B2 net66 VDD pch_mac l=30.0n w=0.17u 
MM4 ZN B3 net65 VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN B3 net65 VDD pch_mac l=30.0n w=0.17u 
MM4_3 ZN B3 net65 VDD pch_mac l=30.0n w=0.17u 
MM4_4 ZN B3 net65 VDD pch_mac l=30.0n w=0.17u 
MM6 net66 B1 net69 VDD pch_mac l=30.0n w=0.17u 
MM6_2 net66 B1 net69 VDD pch_mac l=30.0n w=0.17u 
MM6_3 net66 B1 net69 VDD pch_mac l=30.0n w=0.17u 
MM6_4 net66 B1 net69 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT INVD2 I ZN VDD VSS
MM1 ZN I VSS VSS nch_mac l=30.0n w=0.14u 
MM1_2 ZN I VSS VSS nch_mac l=30.0n w=0.14u 
MM0 ZN I VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 ZN I VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT IOA21D2 A1 A2 B ZN VDD VSS
MM8 net040 net28 VSS VSS nch_mac l=30.0n w=0.14u
MM9 ZN B net040 VSS nch_mac l=30.0n w=0.14u
MM0 net28 A1 net51 VSS nch_mac l=30.0n w=0.14u
MM1 net51 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM6 net39 net28 VSS VSS nch_mac l=30.0n w=0.14u
MM7 ZN B net39 VSS nch_mac l=30.0n w=0.14u
MM5 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM5_2 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM4 ZN net28 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN net28 VDD VDD pch_mac l=30.0n w=0.17u 
MM2 net28 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM3 net28 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT IOA22D2 A1 A2 B1 B2 ZN VDD VSS
MM9 net66 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 net66 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 ZN net30 net66 VSS nch_mac l=30.0n w=0.14u 
MM7_2 ZN net30 net66 VSS nch_mac l=30.0n w=0.14u 
MM6 net66 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 net66 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net30 A2 net50 VSS nch_mac l=30.0n w=0.14u
MM1 net50 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM10 net060 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM11 ZN B2 net060 VDD pch_mac l=30.0n w=0.17u
MM4 net46 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM5 ZN B2 net46 VDD pch_mac l=30.0n w=0.17u
MM8 ZN net30 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_2 ZN net30 VDD VDD pch_mac l=30.0n w=0.17u 
MM2 net30 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM3 net30 A1 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LHCNDD2 D E CDN Q QN VDD VSS
MM25 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM23 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM23_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM22 Q net82 VSS VSS nch_mac l=30.0n w=0.14u 
MM22_2 Q net82 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net150 VSS nch_mac l=30.0n w=0.155u
MM5 net150 D net146 VSS nch_mac l=30.0n w=0.155u
MM7 net146 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM11 net82 qf VSS VSS nch_mac l=30.0n w=140.0n
MM18 qf_x clkb net125 VSS nch_mac l=30.0n w=0.12u
MM19 net118 qf net125 VSS nch_mac l=30.0n w=0.12u
MM20 net118 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM26 clkb E VDD VDD pch_mac l=30.0n w=0.17u
MM24 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM24_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM21 Q net82 VDD VDD pch_mac l=30.0n w=0.17u 
MM21_2 Q net82 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net97 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkb net97 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM10 net82 qf VDD VDD pch_mac l=30.0n w=0.17u
MM16 VDD qf net69 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkbb net69 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT LHCNDQD2 D E CDN Q VDD VSS
MM25 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM20 net92 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM19 net92 qf net91 VSS nch_mac l=30.0n w=0.12u
MM18 qf_x clkb net91 VSS nch_mac l=30.0n w=0.12u
MM12 Q net80 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net80 VSS VSS nch_mac l=30.0n w=0.14u 
MM11 net80 qf VSS VSS nch_mac l=30.0n w=140.0n
MM9 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM7 net71 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM5 net68 D net71 VSS nch_mac l=30.0n w=0.155u
MM4 qf_x clkbb net68 VSS nch_mac l=30.0n w=0.155u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM26 clkb E VDD VDD pch_mac l=30.0n w=0.17u
MM17 qf_x clkbb net139 VDD pch_mac l=30.0n w=0.12u
MM16 VDD qf net139 VDD pch_mac l=30.0n w=0.12u
MM13 Q net80 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net80 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 net80 qf VDD VDD pch_mac l=30.0n w=0.17u
MM8 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkb net112 VDD pch_mac l=30.0n w=0.25u
MM2 net112 D VDD VDD pch_mac l=30.0n w=0.25u
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LHCSNDD2 D E CDN SDN Q QN VDD VSS
MM27 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM26 net0126 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net0106 VSS nch_mac l=30.0n w=0.155u
MM5 net0106 D net0102 VSS nch_mac l=30.0n w=0.155u
MM7 net0102 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net0126 VSS nch_mac l=30.0n w=0.14u
MM11 net0150 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net0150 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net0150 VSS VSS nch_mac l=30.0n w=0.14u 
MM15 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkb net081 VSS nch_mac l=30.0n w=0.12u
MM19 net074 qf net081 VSS nch_mac l=30.0n w=0.12u
MM20 net074 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM28 clkb E VDD VDD pch_mac l=30.0n w=0.17u
MM25 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net0165 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkb net0165 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net0150 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net0150 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net0150 VDD VDD pch_mac l=30.0n w=0.17u 
MM14 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net0137 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkbb net0137 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT LHCSNDQD2 D E CDN SDN Q VDD VSS
MM27 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM26 net0133 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net0138 VSS nch_mac l=30.0n w=0.155u
MM5 net0138 D net0134 VSS nch_mac l=30.0n w=0.155u
MM7 net0134 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net0133 VSS nch_mac l=30.0n w=0.14u
MM11 net0126 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net0126 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net0126 VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkb net0117 VSS nch_mac l=30.0n w=0.12u
MM19 net0114 qf net0117 VSS nch_mac l=30.0n w=0.12u
MM20 net0114 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM28 clkb E VDD VDD pch_mac l=30.0n w=0.17u
MM25 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net089 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkb net089 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net0126 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net0126 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net0126 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net065 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkbb net065 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT LHD2 D E Q QN VDD VSS
MM9 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM8 qf_x clkb net082 VSS nch_mac l=30.0n w=0.12u
MM0 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net112 VSS nch_mac l=30.0n w=0.155u
MM5 net112 D VSS VSS nch_mac l=30.0n w=0.155u
MM11 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM15 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net082 qf VSS VSS nch_mac l=30.0n w=0.12u
MM17 net050 qf VDD VDD pch_mac l=30.0n w=0.12u
MM2 net80 D VDD VDD pch_mac l=30.0n w=0.26u
MM3 qf_x clkb net80 VDD pch_mac l=30.0n w=0.26u
MM10 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM14 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM7 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM18 qf_x clkbb net050 VDD pch_mac l=30.0n w=0.12u
MM1 clkb E VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LHQD2 D E Q VDD VSS
MM9 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM8 net082 clkb qf_x VSS nch_mac l=30.0n w=0.155u
MM0 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net0201 VSS nch_mac l=30.0n w=0.155u
MM5 net0201 D VSS VSS nch_mac l=30.0n w=0.155u
MM11 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM19 VSS qf net082 VSS nch_mac l=30.0n w=0.155u
MM2 net094 D VDD VDD pch_mac l=30.0n w=0.22u
MM3 qf_x clkb net094 VDD pch_mac l=30.0n w=0.22u
MM10 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net0111 VDD pch_mac l=30.0n w=0.22u
MM7 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM6 net0111 clkbb qf_x VDD pch_mac l=30.0n w=0.22u
MM1 clkb E VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LHQOPTDAD2 D E Q VDD VSS
MM9 net92 EB net090 VSS nch_mac l=30n w=100n
MM12_1 net0123 EP VSS VSS nch_mac l=30n w=210.0n
MM12_2 net0123 EP VSS VSS nch_mac l=30n w=210.0n
MM11 net92 D net0123 VSS nch_mac l=30n w=210.0n
MM7 EP EB VSS VSS nch_mac l=30n w=140.0n
MM10 net0240 net92 VSS VSS nch_mac l=30n w=140.0n
MN11 EB E VSS VSS nch_mac l=30n w=140.0n
MM8 net090 net0240 VSS VSS nch_mac l=30n w=100n
MM13_1 Q net92 VSS VSS nch_mac l=30n w=140.0n
MM13_2 Q net92 VSS VSS nch_mac l=30n w=140.0n
MM0 net92 D net0199 VDD pch_mac l=30n w=135.0n
MM3 net200 net0240 VDD VDD pch_mac l=30n w=100n
MM1 net0240 net92 VDD VDD pch_mac l=30n w=170.0n
MM2_1 Q net92 VDD VDD pch_mac l=30n w=170.0n
MM2_2 Q net92 VDD VDD pch_mac l=30n w=170.0n
MM6 EP EB VDD VDD pch_mac l=30n w=170.0n
MM5 EB E VDD VDD pch_mac l=30n w=170.0n
MP12_1 net0199 EB VDD VDD pch_mac l=30n w=135.0n
MP12_2 net0199 EB VDD VDD pch_mac l=30n w=135.0n
MM4 net92 EP net200 VDD pch_mac l=30n w=100n
.ENDS
.SUBCKT LHSNDD2 D E SDN Q QN VDD VSS
MM7 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM26 net134 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net122 VSS nch_mac l=30.0n w=0.155u
MM5 net122 D VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net134 VSS nch_mac l=30.0n w=0.14u
MM11 net70 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net70 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net70 VSS VSS nch_mac l=30.0n w=0.14u 
MM15 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkb net101 VSS nch_mac l=30.0n w=0.12u
MM19 VSS qf net101 VSS nch_mac l=30.0n w=0.12u
MM6 clkb E VDD VDD pch_mac l=30.0n w=0.17u
MM25 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net81 D VDD VDD pch_mac l=30.0n w=0.26u
MM3 qf_x clkb net81 VDD pch_mac l=30.0n w=0.26u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net70 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net70 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net70 VDD VDD pch_mac l=30.0n w=0.17u 
MM14 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net57 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkbb net57 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT LHSNDQD2 D E SDN Q VDD VSS
MM7 clkb E VSS VSS nch_mac l=30.0n w=0.14u
MM26 net065 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkbb net066 VSS nch_mac l=30.0n w=0.155u
MM5 net066 D VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net065 VSS nch_mac l=30.0n w=0.14u
MM11 net058 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net058 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net058 VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkb net049 VSS nch_mac l=30.0n w=0.12u
MM19 VSS qf net049 VSS nch_mac l=30.0n w=0.12u
MM6 clkb E VDD VDD pch_mac l=30.0n w=0.17u
MM25 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net0110 D VDD VDD pch_mac l=30.0n w=0.26u
MM3 qf_x clkb net0110 VDD pch_mac l=30.0n w=0.26u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net058 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net058 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net058 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net093 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkbb net093 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT LNCNDD2 D EN CDN Q QN VDD VSS
MM21 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net95 VSS nch_mac l=30.0n w=0.155u
MM5 net95 D net91 VSS nch_mac l=30.0n w=0.155u
MM7 net91 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM11 net127 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net127 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net127 VSS VSS nch_mac l=30.0n w=0.14u 
MM15 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkbb net70 VSS nch_mac l=30.0n w=0.12u
MM19 net63 qf net70 VSS nch_mac l=30.0n w=0.12u
MM20 net63 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net142 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkbb net142 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM10 net127 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net127 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net127 VDD VDD pch_mac l=30.0n w=0.17u 
MM14 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net118 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkb net118 VDD pch_mac l=30.0n w=0.12u
MM22 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LNCNDQD2 D EN CDN Q VDD VSS
MM21 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net0117 VSS nch_mac l=30.0n w=0.155u
MM5 net0117 D net0113 VSS nch_mac l=30.0n w=0.155u
MM7 net0113 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM11 net0120 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net0120 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net0120 VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkbb net096 VSS nch_mac l=30.0n w=0.12u
MM19 net089 qf net096 VSS nch_mac l=30.0n w=0.12u
MM20 net089 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net080 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkbb net080 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM10 net0120 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net0120 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net0120 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net056 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkb net056 VDD pch_mac l=30.0n w=0.12u
MM22 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LNCSNDD2 D EN CDN SDN Q QN VDD VSS
MM28 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM26 net118 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM23 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM23_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM22 Q net150 VSS VSS nch_mac l=30.0n w=0.14u 
MM22_2 Q net150 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net138 VSS nch_mac l=30.0n w=0.155u
MM5 net138 D net142 VSS nch_mac l=30.0n w=0.155u
MM7 net142 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net118 VSS nch_mac l=30.0n w=0.14u
MM11 net150 qf VSS VSS nch_mac l=30.0n w=140.0n
MM18 qf_x clkbb net169 VSS nch_mac l=30.0n w=0.12u
MM19 net170 qf net169 VSS nch_mac l=30.0n w=0.12u
MM20 net170 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM25 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM24 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM24_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM21 Q net150 VDD VDD pch_mac l=30.0n w=0.17u 
MM21_2 Q net150 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net81 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkbb net81 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net150 qf VDD VDD pch_mac l=30.0n w=0.17u
MM16 VDD qf net109 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkb net109 VDD pch_mac l=30.0n w=0.12u
MM27 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LNCSNDQD2 D EN CDN SDN Q VDD VSS
MM28 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM26 net76 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net81 VSS nch_mac l=30.0n w=0.155u
MM5 net81 D net77 VSS nch_mac l=30.0n w=0.155u
MM7 net77 CDN VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net76 VSS nch_mac l=30.0n w=0.14u
MM11 net121 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net121 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net121 VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkbb net60 VSS nch_mac l=30.0n w=0.12u
MM19 net53 qf net60 VSS nch_mac l=30.0n w=0.12u
MM20 net53 CDN VSS VSS nch_mac l=30.0n w=0.12u
MM25 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net136 D VDD VDD pch_mac l=30.0n w=0.25u
MM3 qf_x clkbb net136 VDD pch_mac l=30.0n w=0.25u
MM6 qf_x CDN VDD VDD pch_mac l=30.0n w=0.25u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net121 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net121 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net121 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 VDD qf net112 VDD pch_mac l=30.0n w=0.12u
MM17 qf_x clkb net112 VDD pch_mac l=30.0n w=0.12u
MM27 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LND2 D EN Q QN VDD VSS
MM6 net77 qf VSS VSS nch_mac l=30.0n w=0.12u
MM8 qf_x clkbb net77 VSS nch_mac l=30.0n w=0.12u
MM9 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net58 VSS nch_mac l=30.0n w=0.155u
MM5 net58 D VSS VSS nch_mac l=30.0n w=0.155u
MM11 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM15 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkb net110 VDD pch_mac l=30.0n w=0.12u
MM17 net110 qf VDD VDD pch_mac l=30.0n w=0.12u
MM2 net120 D VDD VDD pch_mac l=30.0n w=0.26u
MM3 qf_x clkbb net120 VDD pch_mac l=30.0n w=0.26u
MM10 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM14 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM7 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM1 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LNQD2 D EN Q VDD VSS
MM6 net70 qf VSS VSS nch_mac l=30.0n w=0.155u
MM8 qf_x clkbb net70 VSS nch_mac l=30.0n w=0.155u
MM9 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net90 VSS nch_mac l=30.0n w=0.155u
MM5 net90 D VSS VSS nch_mac l=30.0n w=0.155u
MM11 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkb net42 VDD pch_mac l=30.0n w=0.22u
MM17 net42 qf VDD VDD pch_mac l=30.0n w=0.22u
MM2 net53 D VDD VDD pch_mac l=30.0n w=0.22u
MM3 qf_x clkbb net53 VDD pch_mac l=30.0n w=0.22u
MM10 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM7 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM1 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LNSNDD2 D EN SDN Q QN VDD VSS
MM15 net128 qf VSS VSS nch_mac l=30.0n w=0.12u
MM22 net116 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net109 VSS nch_mac l=30.0n w=0.155u
MM5 net109 D VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net116 VSS nch_mac l=30.0n w=0.14u
MM11 net73 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net73 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net73 VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkbb net128 VSS nch_mac l=30.0n w=0.12u
MM7 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM19 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM16 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
MM21 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net61 D VDD VDD pch_mac l=30.0n w=0.26u
MM3 qf_x clkbb net61 VDD pch_mac l=30.0n w=0.26u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net73 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net73 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net73 VDD VDD pch_mac l=30.0n w=0.17u 
MM17 qf_x clkb net85 VDD pch_mac l=30.0n w=0.12u
MM14 net85 qf VDD VDD pch_mac l=30.0n w=0.12u
MM6 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT LNSNDQD2 D EN SDN Q VDD VSS
MM15 net052 qf VSS VSS nch_mac l=30.0n w=0.12u
MM22 net064 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM4 qf_x clkb net065 VSS nch_mac l=30.0n w=0.155u
MM5 net065 D VSS VSS nch_mac l=30.0n w=0.155u
MM9 qf SDN net064 VSS nch_mac l=30.0n w=0.14u
MM11 net057 qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 Q net057 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 Q net057 VSS VSS nch_mac l=30.0n w=0.14u 
MM18 qf_x clkbb net052 VSS nch_mac l=30.0n w=0.12u
MM19 clkb EN VSS VSS nch_mac l=30.0n w=0.14u
MM16 clkb EN VDD VDD pch_mac l=30.0n w=0.17u
MM21 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM1 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM2 net0108 D VDD VDD pch_mac l=30.0n w=0.26u
MM3 qf_x clkbb net0108 VDD pch_mac l=30.0n w=0.26u
MM8 qf SDN VDD VDD pch_mac l=30.0n w=0.17u
MM10 net057 qf VDD VDD pch_mac l=30.0n w=0.17u
MM13 Q net057 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Q net057 VDD VDD pch_mac l=30.0n w=0.17u 
MM17 qf_x clkb net085 VDD pch_mac l=30.0n w=0.12u
MM14 net085 qf VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT MAOI222D2 A B C ZN VDD VSS
MM4 ZN A net33 VSS nch_mac l=30.0n w=0.14u 
MM4_2 ZN A net33 VSS nch_mac l=30.0n w=0.14u 
MM0 net33 B VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 net33 B VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net41 A ZN VSS nch_mac l=30.0n w=0.14u 
MM6_2 net41 A ZN VSS nch_mac l=30.0n w=0.14u 
MM9 net41 C VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 net41 C VSS VSS nch_mac l=30.0n w=0.14u 
MM8 net41 B ZN VSS nch_mac l=30.0n w=0.14u 
MM8_2 net41 B ZN VSS nch_mac l=30.0n w=0.14u 
MM7 net16 B VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 net16 B VDD VDD pch_mac l=30.0n w=0.17u 
MM1 ZN A net16 VDD pch_mac l=30.0n w=0.17u 
MM1_2 ZN A net16 VDD pch_mac l=30.0n w=0.17u 
MM2 net25 C VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 net25 C VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net25 A ZN VDD pch_mac l=30.0n w=0.17u 
MM3_2 net25 A ZN VDD pch_mac l=30.0n w=0.17u 
MM5 net25 B ZN VDD pch_mac l=30.0n w=0.17u 
MM5_2 net25 B ZN VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT MAOI22D2 A1 A2 B1 B2 ZN VDD VSS
MM10 ZN A1 net044 VSS nch_mac l=30.0n w=0.14u
MM11 net044 A2 VSS VSS nch_mac l=30.0n w=140n
MM6 ZN A1 net24 VSS nch_mac l=30.0n w=0.14u
MM9 net12 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net12 B1 VSS VSS nch_mac l=30.0n w=0.14u
MM4 ZN net12 VSS VSS nch_mac l=30.0n w=0.14u 
MM4_2 ZN net12 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net24 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM1 ZN A2 net31 VDD pch_mac l=30.0n w=0.17u 
MM1_2 ZN A2 net31 VDD pch_mac l=30.0n w=0.17u 
MM7 net47 B2 VDD VDD pch_mac l=30.0n w=0.17u
MM0 ZN A1 net31 VDD pch_mac l=30.0n w=0.17u 
MM0_2 ZN A1 net31 VDD pch_mac l=30.0n w=0.17u 
MM2 net31 net12 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 net31 net12 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net12 B1 net47 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT MOAI22D2 A1 A2 B1 B2 ZN VDD VSS
MM5 net12 B1 net36 VSS nch_mac l=30.0n w=0.14u
MM9 net40 A2 ZN VSS nch_mac l=30.0n w=0.14u 
MM9_2 net40 A2 ZN VSS nch_mac l=30.0n w=0.14u 
MM6 net36 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM3 net40 net12 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 net40 net12 VSS VSS nch_mac l=30.0n w=0.14u 
MM4 net40 A1 ZN VSS nch_mac l=30.0n w=0.14u 
MM4_2 net40 A1 ZN VSS nch_mac l=30.0n w=0.14u 
MM7 net12 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM8 net12 B2 VDD VDD pch_mac l=30.0n w=0.17u
MM0 ZN net12 VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 ZN net12 VDD VDD pch_mac l=30.0n w=0.17u 
MM1 VDD A2 net24 VDD pch_mac l=30.0n w=0.17u 
MM1_2 VDD A2 net24 VDD pch_mac l=30.0n w=0.17u 
MM2 net24 A1 ZN VDD pch_mac l=30.0n w=0.17u 
MM2_2 net24 A1 ZN VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT MUX2D2 I0 I1 S Z VDD VSS
MM58 Z net066 VSS VSS nch_mac l=30.0n w=0.14u 
MM58_2 Z net066 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net43 S VSS VSS nch_mac l=30.0n w=0.22u
MM5 net51 I0 VSS VSS nch_mac l=30.0n w=0.22u
MM13 net55 I1 VSS VSS nch_mac l=30.0n w=0.14u
MM14 net55 S net066 VSS nch_mac l=30.0n w=0.22u
MM17 net51 net43 net066 VSS nch_mac l=30.0n w=0.22u
MM59 Z net066 VDD VDD pch_mac l=30.0n w=0.17u 
MM59_2 Z net066 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 net43 S VDD VDD pch_mac l=30.0n w=0.305u
MM15 net55 net43 net066 VDD pch_mac l=30.0n w=0.17u
MM1 net51 I0 VDD VDD pch_mac l=30.0n w=0.215u
MM12 net55 I1 VDD VDD pch_mac l=30.0n w=0.17u
MM16 net51 S net066 VDD pch_mac l=30.0n w=0.215u
.ENDS
.SUBCKT MUX2ND2 I0 I1 S ZN VDD VSS
MM38 ZN net093 VSS VSS nch_mac l=30.0n w=0.14u 
MM38_2 ZN net093 VSS VSS nch_mac l=30.0n w=0.14u 
MM17 net27 net35 net54 VSS nch_mac l=30.0n w=0.22u
MM14 net55 S net54 VSS nch_mac l=30.0n w=0.22u
MM13 net55 I1 VSS VSS nch_mac l=30.0n w=0.14u
MM19 net093 net54 VSS VSS nch_mac l=30.0n w=140.0n
MM5 net27 I0 VSS VSS nch_mac l=30.0n w=0.22u
MM7 net35 S VSS VSS nch_mac l=30.0n w=0.22u
MM37 ZN net093 VDD VDD pch_mac l=30.0n w=0.17u 
MM37_2 ZN net093 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net27 S net54 VDD pch_mac l=30.0n w=0.215u
MM18 net093 net54 VDD VDD pch_mac l=30.0n w=0.17u
MM12 net55 I1 VDD VDD pch_mac l=30.0n w=0.17u
MM1 net27 I0 VDD VDD pch_mac l=30.0n w=0.215u
MM15 net55 net35 net54 VDD pch_mac l=30.0n w=0.17u
MM6 net35 S VDD VDD pch_mac l=30.0n w=0.305u
.ENDS
.SUBCKT MUX2NOPTD2 I0 I1 S ZN VDD VSS
MM8_1 net15 net31 ZN VDD pch_mac l=30n w=170.0n
MM8_2 net15 net31 ZN VDD pch_mac l=30n w=170.0n
MM6_1 net19 S ZN VDD pch_mac l=30n w=170.0n
MM6_2 net19 S ZN VDD pch_mac l=30n w=170.0n
MM1_1 net19 I0 VDD VDD pch_mac l=30n w=170.0n
MM1_2 net19 I0 VDD VDD pch_mac l=30n w=170.0n
MM13 net31 S VDD VDD pch_mac l=30n w=170.0n
MM11_1 net15 I1 VDD VDD pch_mac l=30n w=170.0n
MM11_2 net15 I1 VDD VDD pch_mac l=30n w=170.0n
MM12 net31 S VSS VSS nch_mac l=30n w=140.0n
MM9_1 net15 S ZN VSS nch_mac l=30n w=140.0n
MM9_2 net15 S ZN VSS nch_mac l=30n w=140.0n
MM7_1 net19 net31 ZN VSS nch_mac l=30n w=140.0n
MM7_2 net19 net31 ZN VSS nch_mac l=30n w=140.0n
MM0_1 net19 I0 VSS VSS nch_mac l=30n w=140.0n
MM0_2 net19 I0 VSS VSS nch_mac l=30n w=140.0n
MM10_1 net15 I1 VSS VSS nch_mac l=30n w=140.0n
MM10_2 net15 I1 VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT MUX2OPTD2 I0 I1 S Z VDD VSS
MM0 net33 I0 VSS VSS nch_mac l=30n w=140.0n
MM2 net5 I1 VSS VSS nch_mac l=30n w=140.0n
MM5 net25 S VSS VSS nch_mac l=30n w=140.0n
MM7 net33 net25 net48 VSS nch_mac l=30n w=140.0n
MM9 net5 S net48 VSS nch_mac l=30n w=140.0n
MM11_1 Z net48 VSS VSS nch_mac l=30n w=140.0n
MM11_2 Z net48 VSS VSS nch_mac l=30n w=140.0n
MM1 net33 I0 VDD VDD pch_mac l=30n w=310.0n
MM3 net5 I1 VDD VDD pch_mac l=30n w=170.0n
MM4 net25 S VDD VDD pch_mac l=30n w=170.0n
MM6 net33 S net48 VDD pch_mac l=30n w=310.0n
MM8 net5 net25 net48 VDD pch_mac l=30n w=310.0n
MM10_1 Z net48 VDD VDD pch_mac l=30n w=170.0n
MM10_2 Z net48 VDD VDD pch_mac l=30n w=170.0n
.ENDS
.SUBCKT MUX3D2 I0 I1 I2 S0 S1 Z VDD VSS
MM24 Z net087 VSS VSS nch_mac l=30.0n w=0.14u 
MM24_2 Z net087 VSS VSS nch_mac l=30.0n w=0.14u 
MM20 net61 S1 VSS VSS nch_mac l=30.0n w=0.14u
MM0 net21 I2 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net48 net61 net087 VSS nch_mac l=30.0n w=0.14u
MM8 net21 S1 net087 VSS nch_mac l=30.0n w=140.0n
MM7 net33 S0 VSS VSS nch_mac l=30.0n w=0.14u
MM5 net85 I0 VSS VSS nch_mac l=30.0n w=0.21u
MM13 net89 I1 VSS VSS nch_mac l=30.0n w=0.14u
MM14 net89 S0 net48 VSS nch_mac l=30.0n w=0.14u
MM17 net85 net33 net48 VSS nch_mac l=30.0n w=0.14u
MM25 Z net087 VDD VDD pch_mac l=30.0n w=0.17u 
MM25_2 Z net087 VDD VDD pch_mac l=30.0n w=0.17u 
MM21 net61 S1 VDD VDD pch_mac l=30.0n w=0.17u
MM2 net21 I2 VDD VDD pch_mac l=30.0n w=0.17u
MM11 net48 S1 net087 VDD pch_mac l=30.0n w=0.17u
MM10 net21 net61 net087 VDD pch_mac l=30.0n w=0.17u
MM6 net33 S0 VDD VDD pch_mac l=30.0n w=0.17u
MM15 net89 net33 net48 VDD pch_mac l=30.0n w=0.17u
MM1 net85 I0 VDD VDD pch_mac l=30.0n w=0.17u
MM12 net89 I1 VDD VDD pch_mac l=30.0n w=0.17u
MM16 net85 S0 net48 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT MUX3ND2 I0 I1 I2 S0 S1 ZN VDD VSS
MM24 ZN net0157 VSS VSS nch_mac l=30.0n w=0.14u 
MM24_2 ZN net0157 VSS VSS nch_mac l=30.0n w=0.14u 
MM17 net77 net33 net72 VSS nch_mac l=30.0n w=0.14u
MM14 net73 S0 net72 VSS nch_mac l=30.0n w=0.14u
MM13 net73 I1 VSS VSS nch_mac l=30.0n w=0.14u
MM5 net77 I0 VSS VSS nch_mac l=30.0n w=0.21u
MM7 net33 S0 VSS VSS nch_mac l=30.0n w=0.14u
MM0 net85 I2 VSS VSS nch_mac l=30.0n w=0.14u
MM20 net89 S1 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net85 S1 net96 VSS nch_mac l=30.0n w=140.0n
MM9 net72 net89 net96 VSS nch_mac l=30.0n w=0.14u
MM4 net0157 net96 VSS VSS nch_mac l=30.0n w=0.14u
MM25 ZN net0157 VDD VDD pch_mac l=30.0n w=0.17u 
MM25_2 ZN net0157 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net77 S0 net72 VDD pch_mac l=30.0n w=0.17u
MM12 net73 I1 VDD VDD pch_mac l=30.0n w=0.17u
MM1 net77 I0 VDD VDD pch_mac l=30.0n w=0.17u
MM15 net73 net33 net72 VDD pch_mac l=30.0n w=0.17u
MM6 net33 S0 VDD VDD pch_mac l=30.0n w=0.17u
MM2 net85 I2 VDD VDD pch_mac l=30.0n w=0.17u
MM21 net89 S1 VDD VDD pch_mac l=30.0n w=0.17u
MM10 net85 net89 net96 VDD pch_mac l=30.0n w=0.17u
MM11 net72 S1 net96 VDD pch_mac l=30.0n w=0.17u
MM19 net0157 net96 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT MUX4D2 I0 I1 I2 I3 S0 S1 Z VDD VSS
MM3 Z net0178 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 Z net0178 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net94 I1 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 net94 I1 VSS VSS nch_mac l=30.0n w=0.14u 
MM26 net10 S0 VSS VSS nch_mac l=30.0n w=0.14u
MM10 net70 I3 VSS VSS nch_mac l=30.0n w=0.14u 
MM10_2 net70 I3 VSS VSS nch_mac l=30.0n w=0.14u 
MM9 net66 I2 VSS VSS nch_mac l=30.0n w=0.22u 
MM9_2 net66 I2 VSS VSS nch_mac l=30.0n w=0.22u 
MM33 net66 net10 net81 VSS nch_mac l=30.0n w=0.14u
MM34 net70 S0 net81 VSS nch_mac l=30.0n w=0.14u
MM38 net30 S1 VSS VSS nch_mac l=30.0n w=0.14u
MM39 net81 S1 net0178 VSS nch_mac l=30.0n w=0.14u
MM40 net109 net30 net0178 VSS nch_mac l=30.0n w=0.14u
MM17 net110 net10 net109 VSS nch_mac l=30.0n w=0.14u
MM14 net94 S0 net109 VSS nch_mac l=30.0n w=0.14u
MM5 net110 I0 VSS VSS nch_mac l=30.0n w=0.22u 
MM5_2 net110 I0 VSS VSS nch_mac l=30.0n w=0.22u 
MM0 Z net0178 VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 Z net0178 VDD VDD pch_mac l=30.0n w=0.17u 
MM25 net10 S0 VDD VDD pch_mac l=30.0n w=0.17u
MM8 net66 I2 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_2 net66 I2 VDD VDD pch_mac l=30.0n w=0.17u 
MM11 net70 I3 VDD VDD pch_mac l=30.0n w=0.17u 
MM11_2 net70 I3 VDD VDD pch_mac l=30.0n w=0.17u 
MM32 net70 net10 net81 VDD pch_mac l=30.0n w=0.17u
MM35 net30 S1 VDD VDD pch_mac l=30.0n w=0.17u
MM36 net81 net30 net0178 VDD pch_mac l=30.0n w=0.155u
MM37 net109 S1 net0178 VDD pch_mac l=30.0n w=0.155u
MM16 net110 S0 net109 VDD pch_mac l=30.0n w=0.17u
MM1 net110 I0 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 net110 I0 VDD VDD pch_mac l=30.0n w=0.17u 
MM15 net94 net10 net109 VDD pch_mac l=30.0n w=0.17u
MM31 net66 S0 net81 VDD pch_mac l=30.0n w=0.17u
MM7 net94 I1 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 net94 I1 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT MUX4ND2 I0 I1 I2 I3 S0 S1 ZN VDD VSS
MM13 ZN net0132 VSS VSS nch_mac l=30.0n w=0.14u 
MM13_2 ZN net0132 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net18 I0 VSS VSS nch_mac l=30.0n w=0.175u
MM14 net30 S0 net25 VSS nch_mac l=30.0n w=0.22u
MM17 net18 net126 net25 VSS nch_mac l=30.0n w=0.22u
MM24 net30 I1 VSS VSS nch_mac l=30.0n w=0.22u
MM40 net70 net102 net0132 VSS nch_mac l=30.0n w=0.14u
MM39 net66 S1 net0132 VSS nch_mac l=30.0n w=0.14u
MM38 net102 S1 VSS VSS nch_mac l=30.0n w=0.16u
MM34 net54 S0 net49 VSS nch_mac l=30.0n w=0.14u
MM33 net58 net126 net49 VSS nch_mac l=30.0n w=0.14u
MM30 net54 I3 VSS VSS nch_mac l=30.0n w=140.0n
MM28 net58 I2 VSS VSS nch_mac l=30.0n w=0.16u
MM26 net126 S0 VSS VSS nch_mac l=30.0n w=0.14u
MM4 net66 net49 VSS VSS nch_mac l=30.0n w=0.14u
MM2 net70 net25 VSS VSS nch_mac l=30.0n w=0.14u
MM12 ZN net0132 VDD VDD pch_mac l=30.0n w=0.17u 
MM12_2 ZN net0132 VDD VDD pch_mac l=30.0n w=0.17u 
MM15 net30 net126 net25 VDD pch_mac l=30.0n w=0.285u
MM1 net18 I0 VDD VDD pch_mac l=30.0n w=0.175u
MM16 net18 S0 net25 VDD pch_mac l=30.0n w=0.175u
MM37 net70 S1 net0132 VDD pch_mac l=30.0n w=0.17u
MM36 net66 net102 net0132 VDD pch_mac l=30.0n w=170.0n
MM35 net102 S1 VDD VDD pch_mac l=30.0n w=0.17u
MM31 net58 S0 net49 VDD pch_mac l=30.0n w=0.175u
MM23 net30 I1 VDD VDD pch_mac l=30.0n w=0.295u
MM32 net54 net126 net49 VDD pch_mac l=30.0n w=0.22u
MM27 net58 I2 VDD VDD pch_mac l=30.0n w=0.175u
MM29 net54 I3 VDD VDD pch_mac l=30.0n w=0.17u
MM25 net126 S0 VDD VDD pch_mac l=30.0n w=0.175u
MM0 net70 net25 VDD VDD pch_mac l=30.0n w=170.0n
MM3 net66 net49 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT ND2D2 A1 A2 ZN VDD VSS
MM4 ZN A1 net026 VSS nch_mac l=30.0n w=0.14u 
MM4_2 ZN A1 net026 VSS nch_mac l=30.0n w=0.14u 
MM9 net026 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 net026 A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM1 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM2 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT ND2OPTIBD2 A1 A2 ZN VDD VSS
MM9_1 net026 A2 VSS VSS nch_mac l=30n w=140.0n
MM9_2 net026 A2 VSS VSS nch_mac l=30n w=140.0n
MM4_1 ZN A1 net026 VSS nch_mac l=30n w=140.0n
MM4_2 ZN A1 net026 VSS nch_mac l=30n w=140.0n
MM2_1 ZN A2 VDD VDD pch_mac l=30n w=240.0n
MM2_2 ZN A2 VDD VDD pch_mac l=30n w=240.0n
MM1_1 ZN A1 VDD VDD pch_mac l=30n w=240.0n
MM1_2 ZN A1 VDD VDD pch_mac l=30n w=240.0n
.ENDS
.SUBCKT ND2OPTPAD2 A1 A2 ZN VDD VSS
MM7_1 net045 A2 VSS VSS nch_mac l=30n w=140.0n
MM7_2 net045 A2 VSS VSS nch_mac l=30n w=140.0n
MM7_3 net045 A2 VSS VSS nch_mac l=30n w=140.0n
MM7_4 net045 A2 VSS VSS nch_mac l=30n w=140.0n
MM7_5 net045 A2 VSS VSS nch_mac l=30n w=140.0n
MM7_6 net045 A2 VSS VSS nch_mac l=30n w=140.0n
MM10_1 ZN A1 net045 VSS nch_mac l=30n w=140.0n
MM10_2 ZN A1 net045 VSS nch_mac l=30n w=140.0n
MM1_1 ZN A1 VDD VDD pch_mac l=30n w=170.0n
MM1_2 ZN A1 VDD VDD pch_mac l=30n w=170.0n
MM8_1 ZN A2 VDD VDD pch_mac l=30n w=170.0n
MM8_2 ZN A2 VDD VDD pch_mac l=30n w=170.0n
.ENDS
.SUBCKT ND3D2 A1 A2 A3 ZN VDD VSS
MM18 net031 A2 net023 VSS nch_mac l=30.0n w=140.0n
MM19 ZN A1 net031 VSS nch_mac l=30.0n w=140.0n
MM20 net023 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM15 net40 A2 net32 VSS nch_mac l=30.0n w=0.14u
MM16 ZN A1 net40 VSS nch_mac l=30.0n w=0.14u
MM17 net32 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM9 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_2 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM14 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM14_2 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 ZN A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 ZN A3 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT ND3OPTPAD2 A1 A2 A3 ZN VDD VSS
MM2_1 net041 A3 VSS VSS nch_mac l=30n w=140.0n
MM2_2 net041 A3 VSS VSS nch_mac l=30n w=140.0n
MM2_3 net041 A3 VSS VSS nch_mac l=30n w=140.0n
MM2_4 net041 A3 VSS VSS nch_mac l=30n w=140.0n
MM7_1 net045 A2 net041 VSS nch_mac l=30n w=140.0n
MM7_2 net045 A2 net041 VSS nch_mac l=30n w=140.0n
MM7_3 net045 A2 net041 VSS nch_mac l=30n w=140.0n
MM7_4 net045 A2 net041 VSS nch_mac l=30n w=140.0n
MM10_1 ZN A1 net045 VSS nch_mac l=30n w=140.0n
MM10_2 ZN A1 net045 VSS nch_mac l=30n w=140.0n
MM1_1 ZN A1 VDD VDD pch_mac l=30n w=170.0n
MM1_2 ZN A1 VDD VDD pch_mac l=30n w=170.0n
MM8_1 ZN A2 VDD VDD pch_mac l=30n w=170.0n
MM8_2 ZN A2 VDD VDD pch_mac l=30n w=170.0n
MM19_1 ZN A3 VDD VDD pch_mac l=30n w=170.0n
MM19_2 ZN A3 VDD VDD pch_mac l=30n w=170.0n
.ENDS
.SUBCKT ND4D2 A1 A2 A3 A4 ZN VDD VSS
MM9 net123 A4 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 net123 A4 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net119 A3 net123 VSS nch_mac l=30.0n w=0.14u 
MM7_2 net119 A3 net123 VSS nch_mac l=30.0n w=0.14u 
MM22 ZN A1 net111 VSS nch_mac l=30.0n w=0.14u 
MM22_2 ZN A1 net111 VSS nch_mac l=30.0n w=0.14u 
MM23 net111 A2 net119 VSS nch_mac l=30.0n w=0.14u 
MM23_2 net111 A2 net119 VSS nch_mac l=30.0n w=0.14u 
MM8 ZN A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM8_2 ZN A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM10_2 ZN A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM11 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM11_2 ZN A1 VDD VDD pch_mac l=30.0n w=0.17u 
MM12 ZN A4 VDD VDD pch_mac l=30.0n w=0.17u 
MM12_2 ZN A4 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT NR2D2 A1 A2 ZN VDD VSS
MM18 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM18_2 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM19 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM19_2 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 ZN A1 net034 VDD pch_mac l=30.0n w=0.17u 
MM5_2 ZN A1 net034 VDD pch_mac l=30.0n w=0.17u 
MM6 net034 A2 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 net034 A2 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT NR2OPTIBD2 A1 A2 ZN VDD VSS
MM19_1 ZN A1 VSS VSS nch_mac l=30n w=240.0n
MM19_2 ZN A1 VSS VSS nch_mac l=30n w=240.0n
MM18_1 ZN A2 VSS VSS nch_mac l=30n w=240.0n
MM18_2 ZN A2 VSS VSS nch_mac l=30n w=240.0n
MM17 net034 A2 VDD VDD pch_mac l=30n w=170.0n
MM6 net034 A2 VDD VDD pch_mac l=30n w=170.0n
MM16 ZN A1 net034 VDD pch_mac l=30n w=170.0n
MM5 ZN A1 net034 VDD pch_mac l=30n w=170.0n
.ENDS
.SUBCKT NR2OPTPAD2 A1 A2 ZN VDD VSS
MM2_1 ZN A1 VSS VSS nch_mac l=30n w=140.0n
MM2_2 ZN A1 VSS VSS nch_mac l=30n w=140.0n
MM7_1 ZN A2 VSS VSS nch_mac l=30n w=140.0n
MM7_2 ZN A2 VSS VSS nch_mac l=30n w=140.0n
MM1_1 net040 A2 VDD VDD pch_mac l=30n w=170.0n
MM1_2 net040 A2 VDD VDD pch_mac l=30n w=170.0n
MM8 ZN A1 net040 VDD pch_mac l=30n w=170.0n
MM20_1 net021 A2 VDD VDD pch_mac l=30n w=170.0n
MM20_2 net021 A2 VDD VDD pch_mac l=30n w=170.0n
MM19 ZN A1 net021 VDD pch_mac l=30n w=170.0n
.ENDS
.SUBCKT NR3D2 A1 A2 A3 ZN VDD VSS
MM12 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM13 ZN A3 VSS VSS nch_mac l=30.0n w=0.14u 
MM13_2 ZN A3 VSS VSS nch_mac l=30.0n w=0.14u 
MM14 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM14_2 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM3 net78 A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_2 net78 A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_3 net78 A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM3_4 net78 A3 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 ZN A1 net82 VDD pch_mac l=30.0n w=0.17u 
MM10_2 ZN A1 net82 VDD pch_mac l=30.0n w=0.17u 
MM10_3 ZN A1 net82 VDD pch_mac l=30.0n w=0.17u 
MM10_4 ZN A1 net82 VDD pch_mac l=30.0n w=0.17u 
MM11 net82 A2 net78 VDD pch_mac l=30.0n w=0.17u 
MM11_2 net82 A2 net78 VDD pch_mac l=30.0n w=0.17u 
MM11_3 net82 A2 net78 VDD pch_mac l=30.0n w=0.17u 
MM11_4 net82 A2 net78 VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT NR3OPTPAD2 A1 A2 A3 ZN VDD VSS
MM2_1 ZN A3 VSS VSS nch_mac l=30n w=140.0n
MM2_2 ZN A3 VSS VSS nch_mac l=30n w=140.0n
MM7_1 ZN A1 VSS VSS nch_mac l=30n w=140.0n
MM7_2 ZN A1 VSS VSS nch_mac l=30n w=140.0n
MM10_1 ZN A2 VSS VSS nch_mac l=30n w=140.0n
MM10_2 ZN A2 VSS VSS nch_mac l=30n w=140.0n
MM1_1 net040 A3 VDD VDD pch_mac l=30n w=170.0n
MM1_2 net040 A3 VDD VDD pch_mac l=30n w=170.0n
MM1_3 net040 A3 VDD VDD pch_mac l=30n w=170.0n
MM1_4 net040 A3 VDD VDD pch_mac l=30n w=170.0n
MM1_5 net040 A3 VDD VDD pch_mac l=30n w=170.0n
MM8_1 net025 A2 net040 VDD pch_mac l=30n w=170.0n
MM8_2 net025 A2 net040 VDD pch_mac l=30n w=170.0n
MM8_3 net025 A2 net040 VDD pch_mac l=30n w=170.0n
MM8_4 net025 A2 net040 VDD pch_mac l=30n w=170.0n
MM19_1 ZN A1 net025 VDD pch_mac l=30n w=170.0n
MM19_2 ZN A1 net025 VDD pch_mac l=30n w=170.0n
.ENDS
.SUBCKT NR4D2 A1 A2 A3 A4 ZN VDD VSS
MM2 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A1 VSS VSS nch_mac l=30.0n w=0.14u 
MM9 ZN A3 VSS VSS nch_mac l=30.0n w=0.14u 
MM9_2 ZN A3 VSS VSS nch_mac l=30.0n w=0.14u 
MM8 ZN A4 VSS VSS nch_mac l=30.0n w=0.14u 
MM8_2 ZN A4 VSS VSS nch_mac l=30.0n w=0.14u 
MM1 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM1_2 ZN A2 VSS VSS nch_mac l=30.0n w=0.14u 
MM4 ZN A1 net11 VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN A1 net11 VDD pch_mac l=30.0n w=0.17u 
MM4_3 ZN A1 net11 VDD pch_mac l=30.0n w=0.17u 
MM4_4 ZN A1 net11 VDD pch_mac l=30.0n w=0.17u 
MM7 net19 A3 net15 VDD pch_mac l=30.0n w=0.17u 
MM7_2 net19 A3 net15 VDD pch_mac l=30.0n w=0.17u 
MM7_3 net19 A3 net15 VDD pch_mac l=30.0n w=0.17u 
MM7_4 net19 A3 net15 VDD pch_mac l=30.0n w=0.17u 
MM3 net11 A2 net19 VDD pch_mac l=30.0n w=0.17u 
MM3_2 net11 A2 net19 VDD pch_mac l=30.0n w=0.17u 
MM3_3 net11 A2 net19 VDD pch_mac l=30.0n w=0.17u 
MM3_4 net11 A2 net19 VDD pch_mac l=30.0n w=0.17u 
MM0 net15 A4 VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 net15 A4 VDD VDD pch_mac l=30.0n w=0.17u 
MM0_3 net15 A4 VDD VDD pch_mac l=30.0n w=0.17u 
MM0_4 net15 A4 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT OA211D2 A1 A2 B C Z VDD VSS
MM5 Z net20 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net20 VSS VSS nch_mac l=30.0n w=0.14u 
MM13 net12 C VSS VSS nch_mac l=30.0n w=0.14u
MM12 net23 B net12 VSS nch_mac l=30.0n w=0.14u
MM8 net20 A1 net23 VSS nch_mac l=30.0n w=0.14u
MM9 net20 A2 net23 VSS nch_mac l=30.0n w=0.14u
MM4 Z net20 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net20 VDD VDD pch_mac l=30.0n w=0.17u 
MM10 net20 C VDD VDD pch_mac l=30.0n w=0.17u
MM11 net20 B VDD VDD pch_mac l=30.0n w=0.17u
MM6 net47 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM7 net20 A2 net47 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OA21D2 A1 A2 B Z VDD VSS
MM6 Z net15 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 Z net15 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net18 B VSS VSS nch_mac l=30.0n w=0.14u
MM8 net15 A2 net18 VSS nch_mac l=30.0n w=0.14u
MM9 net15 A1 net18 VSS nch_mac l=30.0n w=0.14u
MM10 Z net15 VDD VDD pch_mac l=30.0n w=0.17u 
MM10_2 Z net15 VDD VDD pch_mac l=30.0n w=0.17u 
MM11 net15 A1 net30 VDD pch_mac l=30.0n w=0.17u
MM12 net30 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM13 net15 B VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OA22D2 A1 A2 B1 B2 Z VDD VSS
MM5 Z net44 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net44 VSS VSS nch_mac l=30.0n w=0.14u 
MM13 net47 B2 VSS VSS nch_mac l=30.0n w=0.14u
MM12 net47 B1 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net44 A2 net47 VSS nch_mac l=30.0n w=0.14u
MM8 net44 A1 net47 VSS nch_mac l=30.0n w=0.14u
MM4 Z net44 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net44 VDD VDD pch_mac l=30.0n w=0.17u 
MM11 net19 B2 VDD VDD pch_mac l=30.0n w=0.17u
MM10 net44 B1 net19 VDD pch_mac l=30.0n w=0.17u
MM7 net44 A1 net23 VDD pch_mac l=30.0n w=0.17u
MM6 net23 A2 VDD VDD pch_mac l=30.0n w=170.0n
.ENDS
.SUBCKT OAI211D2 A1 A2 B C ZN VDD VSS
MM9 net060 C VSS VSS nch_mac l=30.0n w=0.14u
MM10 net39 B net060 VSS nch_mac l=30.0n w=0.14u
MM7 net24 C VSS VSS nch_mac l=30.0n w=0.14u
MM6 net39 B net24 VSS nch_mac l=30.0n w=0.14u
MM58 ZN A2 net39 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A2 net39 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A1 net39 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A1 net39 VSS nch_mac l=30.0n w=0.14u 
MM3 net032 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM8 ZN A2 net032 VDD pch_mac l=30.0n w=0.17u
MM4 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM5 ZN C VDD VDD pch_mac l=30.0n w=0.17u 
MM5_2 ZN C VDD VDD pch_mac l=30.0n w=0.17u 
MM1 net23 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM0 ZN A2 net23 VDD pch_mac l=30.0n w=170.0n
.ENDS
.SUBCKT OAI211OPTREPBD2 A1 A2 B C ZN VDD VSS
MP11_1 ZN A1 net046 VDD pch_mac l=30n w=170.0n
MP11_2 ZN A1 net046 VDD pch_mac l=30n w=170.0n
MP31_1 ZN B VDD VDD pch_mac l=30n w=170.0n
MP31_2 ZN B VDD VDD pch_mac l=30n w=170.0n
MP21_1 ZN C VDD VDD pch_mac l=30n w=170.0n
MP21_2 ZN C VDD VDD pch_mac l=30n w=170.0n
MP12_1 net046 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_2 net046 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_3 net046 A2 VDD VDD pch_mac l=30n w=170.0n
MP12_4 net046 A2 VDD VDD pch_mac l=30n w=170.0n
MN12_1 ZN B net030 VSS nch_mac l=30n w=140.0n
MN12_2 ZN B net030 VSS nch_mac l=30n w=140.0n
MN11_1 net019 A1 VSS VSS nch_mac l=30n w=140.0n
MN11_2 net019 A1 VSS VSS nch_mac l=30n w=140.0n
MN11_3 net019 A1 VSS VSS nch_mac l=30n w=140.0n
MN11_4 net019 A1 VSS VSS nch_mac l=30n w=140.0n
MN21_1 net019 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_2 net019 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_3 net019 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_4 net019 A2 VSS VSS nch_mac l=30n w=140.0n
MN13_1 net030 C net019 VSS nch_mac l=30n w=140.0n
MN13_2 net030 C net019 VSS nch_mac l=30n w=140.0n
MN13_3 net030 C net019 VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT OAI21D2 A1 A2 B ZN VDD VSS
MM3 net30 B VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 net30 B VSS VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A2 net30 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A2 net30 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A1 net30 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A1 net30 VSS nch_mac l=30.0n w=0.14u 
MM4 ZN A1 net031 VDD pch_mac l=30.0n w=0.17u
MM5 net031 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM59 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM59_2 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM0 ZN A1 net14 VDD pch_mac l=30.0n w=170.0n
MM1 net14 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OAI21OPTREPBD2 A1 A2 B ZN VDD VSS
MP11_1 net036 A2 VDD VDD pch_mac l=30n w=170.0n
MP11_2 net036 A2 VDD VDD pch_mac l=30n w=170.0n
MP11_3 net036 A2 VDD VDD pch_mac l=30n w=170.0n
MP11_4 net036 A2 VDD VDD pch_mac l=30n w=170.0n
MP31_1 ZN B VDD VDD pch_mac l=30n w=170.0n
MP31_2 ZN B VDD VDD pch_mac l=30n w=170.0n
MP12_1 ZN A1 net036 VDD pch_mac l=30n w=170.0n
MP12_2 ZN A1 net036 VDD pch_mac l=30n w=170.0n
MN12_1 ZN B net021 VSS nch_mac l=30n w=140.0n
MN12_2 ZN B net021 VSS nch_mac l=30n w=140.0n
MN11_1 net021 A1 VSS VSS nch_mac l=30n w=140.0n
MN11_2 net021 A1 VSS VSS nch_mac l=30n w=140.0n
MN11_3 net021 A1 VSS VSS nch_mac l=30n w=140.0n
MN11_4 net021 A1 VSS VSS nch_mac l=30n w=140.0n
MN21_1 net021 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_2 net021 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_3 net021 A2 VSS VSS nch_mac l=30n w=140.0n
MN21_4 net021 A2 VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT OAI221D2 A1 A2 B1 B2 C ZN VDD VSS
MM7 net20 C VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net20 C VSS VSS nch_mac l=30.0n w=0.14u 
MM9 net24 B1 net20 VSS nch_mac l=30.0n w=0.14u 
MM9_2 net24 B1 net20 VSS nch_mac l=30.0n w=0.14u 
MM5 net24 B2 net20 VSS nch_mac l=30.0n w=0.14u 
MM5_2 net24 B2 net20 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A2 net24 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A2 net24 VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A1 net24 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A1 net24 VSS nch_mac l=30.0n w=0.14u 
MM6 ZN A1 net070 VDD pch_mac l=30.0n w=170.0n
MM10 net070 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM11 net058 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM12 ZN B2 net058 VDD pch_mac l=30.0n w=0.17u
MM4 ZN C VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 ZN C VDD VDD pch_mac l=30.0n w=0.17u 
MM8 net40 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM3 ZN B2 net40 VDD pch_mac l=30.0n w=0.17u
MM0 ZN A1 net44 VDD pch_mac l=30.0n w=170.0n
MM1 net44 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OAI222D2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM7 net45 C2 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net45 C2 VSS VSS nch_mac l=30.0n w=0.14u 
MM10 net45 C1 VSS VSS nch_mac l=30.0n w=0.14u 
MM10_2 net45 C1 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net53 B2 net45 VSS nch_mac l=30.0n w=0.14u 
MM5_2 net53 B2 net45 VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A1 net53 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A1 net53 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A2 net53 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A2 net53 VSS nch_mac l=30.0n w=0.14u 
MM9 net53 B1 net45 VSS nch_mac l=30.0n w=0.14u 
MM9_2 net53 B1 net45 VSS nch_mac l=30.0n w=0.14u 
MM11 net058 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM12 ZN A1 net058 VDD pch_mac l=30.0n w=0.17u
MM13 ZN B2 net054 VDD pch_mac l=30.0n w=0.17u
MM14 net054 B1 VDD VDD pch_mac l=30.0n w=170.0n
MM4 ZN C2 net13 VDD pch_mac l=30.0n w=0.17u
MM6 net13 C1 VDD VDD pch_mac l=30.0n w=170.0n
MM1 net25 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM0 ZN A1 net25 VDD pch_mac l=30.0n w=170.0n
MM3 ZN B2 net29 VDD pch_mac l=30.0n w=0.17u
MM8 net29 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM15 ZN C2 net046 VDD pch_mac l=30.0n w=0.17u
MM16 net046 C1 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OAI22D2 A1 A2 B1 B2 ZN VDD VSS
MM7 net19 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net19 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM6 net19 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 net19 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A1 net19 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A1 net19 VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A2 net19 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A2 net19 VSS nch_mac l=30.0n w=0.14u 
MM3 ZN A1 net059 VDD pch_mac l=30.0n w=0.17u
MM8 net059 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM9 ZN B1 net051 VDD pch_mac l=30.0n w=0.17u
MM10 net051 B2 VDD VDD pch_mac l=30.0n w=0.17u
MM4 ZN B1 net27 VDD pch_mac l=30.0n w=0.17u
MM5 net27 B2 VDD VDD pch_mac l=30.0n w=0.17u
MM0 ZN A1 net35 VDD pch_mac l=30.0n w=170.0n
MM1 net35 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OAI22OPTPBD2 A1 A2 B1 B2 ZN VDD VSS
MM1_1 net050 B2 VDD VDD pch_mac l=30n w=170.0n
MM1_2 net050 B2 VDD VDD pch_mac l=30n w=170.0n
MM1_3 net050 B2 VDD VDD pch_mac l=30n w=170.0n
MM1_4 net050 B2 VDD VDD pch_mac l=30n w=170.0n
MM9_1 ZN B1 net050 VDD pch_mac l=30n w=170.0n
MM9_2 ZN B1 net050 VDD pch_mac l=30n w=170.0n
MM3_1 net042 A2 VDD VDD pch_mac l=30n w=170.0n
MM3_2 net042 A2 VDD VDD pch_mac l=30n w=170.0n
MM3_3 net042 A2 VDD VDD pch_mac l=30n w=170.0n
MM3_4 net042 A2 VDD VDD pch_mac l=30n w=170.0n
MM4_1 ZN A1 net042 VDD pch_mac l=30n w=170.0n
MM4_2 ZN A1 net042 VDD pch_mac l=30n w=170.0n
MM28_1 net022 B1 VSS VSS nch_mac l=30n w=140.0n
MM28_2 net022 B1 VSS VSS nch_mac l=30n w=140.0n
MM28_3 net022 B1 VSS VSS nch_mac l=30n w=140.0n
MM28_4 net022 B1 VSS VSS nch_mac l=30n w=140.0n
MM6_1 ZN A1 net022 VSS nch_mac l=30n w=140.0n
MM6_2 ZN A1 net022 VSS nch_mac l=30n w=140.0n
MM5_1 ZN A2 net022 VSS nch_mac l=30n w=140.0n
MM5_2 ZN A2 net022 VSS nch_mac l=30n w=140.0n
MM2_1 net022 B2 VSS VSS nch_mac l=30n w=140.0n
MM2_2 net022 B2 VSS VSS nch_mac l=30n w=140.0n
MM2_3 net022 B2 VSS VSS nch_mac l=30n w=140.0n
MM2_4 net022 B2 VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT OAI31D2 A1 A2 A3 B ZN VDD VSS
MM8 ZN A3 net27 VSS nch_mac l=30.0n w=0.14u 
MM8_2 ZN A3 net27 VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A1 net27 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A1 net27 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A2 net27 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A2 net27 VSS nch_mac l=30.0n w=0.14u 
MM7 net27 B VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net27 B VSS VSS nch_mac l=30.0n w=0.14u 
MM4 net033 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM6 net029 A2 net033 VDD pch_mac l=30.0n w=170.0n
MM9 ZN A3 net029 VDD pch_mac l=30.0n w=0.17u
MM5 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM5_2 ZN B VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net19 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM1 net23 A2 net19 VDD pch_mac l=30.0n w=0.17u
MM0 ZN A3 net23 VDD pch_mac l=30.0n w=170.0n
.ENDS
.SUBCKT OAI32D2 A1 A2 A3 B1 B2 ZN VDD VSS
MM4 net28 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM4_2 net28 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net28 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net28 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A2 net28 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A2 net28 VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A1 net28 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A1 net28 VSS nch_mac l=30.0n w=0.14u 
MM8 ZN A3 net28 VSS nch_mac l=30.0n w=0.14u 
MM8_2 ZN A3 net28 VSS nch_mac l=30.0n w=0.14u 
MM13 ZN B2 net32 VDD pch_mac l=30.0n w=0.17u
MM12 net32 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM11 net44 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM10 net48 A2 net44 VDD pch_mac l=30.0n w=0.17u
MM9 ZN A3 net48 VDD pch_mac l=30.0n w=0.17u
MM6 net56 B1 VDD VDD pch_mac l=30.0n w=170.0n
MM5 ZN B2 net56 VDD pch_mac l=30.0n w=0.17u
MM0 ZN A3 net60 VDD pch_mac l=30.0n w=170.0n
MM1 net60 A2 net64 VDD pch_mac l=30.0n w=0.17u
MM3 net64 A1 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OAI33D2 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM10 net41 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM10_2 net41 B2 VSS VSS nch_mac l=30.0n w=0.14u 
MM8 ZN A3 net41 VSS nch_mac l=30.0n w=0.14u 
MM8_2 ZN A3 net41 VSS nch_mac l=30.0n w=0.14u 
MM58 ZN A1 net41 VSS nch_mac l=30.0n w=0.14u 
MM58_2 ZN A1 net41 VSS nch_mac l=30.0n w=0.14u 
MM2 ZN A2 net41 VSS nch_mac l=30.0n w=0.14u 
MM2_2 ZN A2 net41 VSS nch_mac l=30.0n w=0.14u 
MM4 net41 B3 VSS VSS nch_mac l=30.0n w=0.14u 
MM4_2 net41 B3 VSS VSS nch_mac l=30.0n w=0.14u 
MM7 net41 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM7_2 net41 B1 VSS VSS nch_mac l=30.0n w=0.14u 
MM11 net055 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM12 net051 B2 net055 VDD pch_mac l=30.0n w=0.17u
MM13 ZN B3 net051 VDD pch_mac l=30.0n w=0.17u
MM16 ZN A3 net039 VDD pch_mac l=30.0n w=0.17u
MM14 net043 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM15 net039 A2 net043 VDD pch_mac l=30.0n w=0.17u
MM5 net17 B1 VDD VDD pch_mac l=30.0n w=0.17u
MM6 net21 B2 net17 VDD pch_mac l=30.0n w=170.0n
MM9 ZN B3 net21 VDD pch_mac l=30.0n w=0.17u
MM3 net29 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM1 net33 A2 net29 VDD pch_mac l=30.0n w=0.17u
MM0 ZN A3 net33 VDD pch_mac l=30.0n w=170.0n
.ENDS
.SUBCKT OR2D2 A1 A2 Z VDD VSS
MM0 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u 
MM8 net26 A2 VSS VSS nch_mac l=30.0n w=140.0n
MM9 net26 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM1 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net26 A1 net13 VDD pch_mac l=30.0n w=0.17u
MM7 net13 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OR3D2 A1 A2 A3 Z VDD VSS
MM0 Z net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM4 net11 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM9 net11 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net11 A1 VSS VSS nch_mac l=30.0n w=140.0n
MM1 Z net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net11 VDD VDD pch_mac l=30.0n w=0.17u 
MM2 net11 A3 net30 VDD pch_mac l=30.0n w=0.17u
MM7 net38 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM3 net30 A2 net38 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT OR4D2 A1 A2 A3 A4 Z VDD VSS
MM6 net28 A4 VSS VSS nch_mac l=30.0n w=0.14u
MM0 Z net28 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net28 VSS VSS nch_mac l=30.0n w=0.14u 
MM8 net28 A1 VSS VSS nch_mac l=30.0n w=140.0n
MM9 net28 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM4 net28 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM5 net23 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM1 Z net28 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net28 VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net27 A3 net19 VDD pch_mac l=30.0n w=0.17u
MM7 net19 A2 net23 VDD pch_mac l=30.0n w=0.17u
MM2 net28 A4 net27 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFCNARD2 SI D SE CP CDN Q QN VDD VSS
MM0 net0110 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM1 qf_x qf net0110 VSS nch_mac l=30.0n w=0.14u
MM47 net82 net0237 net13 VSS nch_mac l=30.0n w=0.175u
MM51 net85 SI VSS VSS nch_mac l=30.0n w=100n
MM75 net18 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.15u
MM76 qf_x qf net18 VSS nch_mac l=30.0n w=0.14u
MM46 mq_x clkb net82 VSS nch_mac l=30.0n w=0.165u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140n
MM66 net42 CDN VSS VSS nch_mac l=30.0n w=100n
MM64 mq_x clkbb net54 VSS nch_mac l=30.0n w=100n
MM57 net0237 SE VSS VSS nch_mac l=30.0n w=0.12u
MM65 net54 mq net42 VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM69 QN net66 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net66 VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net66 clkb qf VSS nch_mac l=30.0n w=0.15u
MM48 net13 D VSS VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.15u
MM73 net66 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM52 net82 SE net85 VSS nch_mac l=30.0n w=100n
MM2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM43 net13 D VDD VDD pch_mac l=30.0n w=0.275u
MM79 mq_x clkb net101 VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net66 clkbb qf VDD pch_mac l=30.0n w=0.14u
MM44 net158 SE net13 VDD pch_mac l=30.0n w=0.275u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM61 net101 mq VDD VDD pch_mac l=30.0n w=120n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.17u
MM41 net161 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net101 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM74 net66 qf_x VDD VDD pch_mac l=30.0n w=0.14u
MM58 net0237 SE VDD VDD pch_mac l=30.0n w=0.275u
MM70 QN net66 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net66 VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkbb net158 VDD pch_mac l=30.0n w=0.22u
MM42 net158 net0237 net161 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFCND2 SI D SE CP CDN Q QN VDD VSS
MM0 net0110 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM1 qf_x qf net0110 VSS nch_mac l=30.0n w=0.245u
MM47 net82 net0237 net13 VSS nch_mac l=30.0n w=0.175u
MM51 net85 SI VSS VSS nch_mac l=30.0n w=100n
MM75 net18 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.245u
MM76 qf_x qf net18 VSS nch_mac l=30.0n w=0.245u
MM46 mq_x clkb net82 VSS nch_mac l=30.0n w=0.165u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM66 net42 CDN VSS VSS nch_mac l=30.0n w=100n
MM64 mq_x clkbb net54 VSS nch_mac l=30.0n w=100n
MM57 net0237 SE VSS VSS nch_mac l=30.0n w=0.12u
MM65 net54 mq net42 VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM69 QN net66 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net66 VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net66 clkb qf VSS nch_mac l=30.0n w=0.155u
MM48 net13 D VSS VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.155u
MM73 net66 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM52 net82 SE net85 VSS nch_mac l=30.0n w=100n
MM2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.12u
MM2B qf_x CDN VDD VDD pch_mac l=30.0n w=0.295u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.295u
MM43 net13 D VDD VDD pch_mac l=30.0n w=0.275u
MM79 mq_x clkb net101 VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net66 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM44 net158 SE net13 VDD pch_mac l=30.0n w=0.275u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.295u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.295u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM61 net101 mq VDD VDD pch_mac l=30.0n w=120.0n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.295u
MM41 net161 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net101 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM74 net66 qf_x VDD VDD pch_mac l=30.0n w=0.3u
MM58 net0237 SE VDD VDD pch_mac l=30.0n w=0.275u
MM70 QN net66 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net66 VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkbb net158 VDD pch_mac l=30.0n w=0.22u
MM42 net158 net0237 net161 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFCNOPTBD2 SI D SE CP CDN Q QN VDD VSS
MM66 net0111 CDN VSS VSS nch_mac l=30n w=100n
MM64 ml_ax clkbb net0110 VSS nch_mac l=30n w=100n
MM65 net0110 ml_b net0111 VSS nch_mac l=30n w=100n
MM53 clkb CP VSS VSS nch_mac l=30n w=140.0n
MM55 clkbb clkb VSS VSS nch_mac l=30n w=140.0n
MM47_1 net034 D VSS VSS nch_mac l=30n w=135.0n
MM47_2 net034 D VSS VSS nch_mac l=30n w=135.0n
MM49_1 ml_b ml_ax VSS VSS nch_mac l=30n w=240.00n
MM49_2 ml_b ml_ax VSS VSS nch_mac l=30n w=240.00n
MM51 net0109 SI VSS VSS nch_mac l=30n w=100n
MM57 net027 SE VSS VSS nch_mac l=30n w=135.0n
MM52 net031 SE net0109 VSS nch_mac l=30n w=100n
MM73 net66 qf_x VSS VSS nch_mac l=30n w=140.0n
MSLTn1 qf clkbb ml_b VSS nch_mac l=30n w=155.00n
MM67 net66 clkb qf VSS nch_mac l=30n w=155.00n
MM69_1 QN net66 VSS VSS nch_mac l=30n w=140.0n
MM69_2 QN net66 VSS VSS nch_mac l=30n w=140.0n
MM71_1 Q qf_x VSS VSS nch_mac l=30n w=140.0n
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=140.0n
MM46 ml_ax clkb net031 VSS nch_mac l=30n w=165.00n
MM76 qf_x qf net0112 VSS nch_mac l=30n w=240.00n
MM75 net0112 CDN VSS VSS nch_mac l=30n w=240.00n
MM27_1 net031 net027 net034 VSS nch_mac l=30n w=210.0n
MM27_2 net031 net027 net034 VSS nch_mac l=30n w=210.0n
MM1 qf_x qf net0108 VSS nch_mac l=30n w=240.00n
MM0 net0108 CDN VSS VSS nch_mac l=30n w=240.00n
MM61 net0116 ml_b VDD VDD pch_mac l=30n w=120.0n
MM79 ml_ax clkb net0116 VDD pch_mac l=30n w=120.0n
MM60 net0116 CDN VDD VDD pch_mac l=30n w=120.0n
MM54 clkb CP VDD VDD pch_mac l=30n w=170.0n
MM56 clkbb clkb VDD VDD pch_mac l=30n w=170.0n
MM58 net027 SE VDD VDD pch_mac l=30n w=170.0n
MM70_1 QN net66 VDD VDD pch_mac l=30n w=170.0n
MM70_2 QN net66 VDD VDD pch_mac l=30n w=170.0n
MM74 net66 qf_x VDD VDD pch_mac l=30n w=300n
MM78 qf_x CDN VDD VDD pch_mac l=30n w=170.0n
MM77_1 qf_x qf VDD VDD pch_mac l=30n w=170.0n
MM77_2 qf_x qf VDD VDD pch_mac l=30n w=170.0n
MM68 net66 clkbb qf VDD pch_mac l=30n w=120.0n
MM72_1 Q qf_x VDD VDD pch_mac l=30n w=170.0n
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=170.0n
MSLTp1 qf clkb ml_b VDD pch_mac l=30n w=295.00n
MM17 net034 D VDD VDD pch_mac l=30n w=170.0n
MM44_1 net032 SE net034 VDD pch_mac l=30n w=240.00n
MM44_2 net032 SE net034 VDD pch_mac l=30n w=240.00n
MM41 net0107 SI VDD VDD pch_mac l=30n w=100n
MM42 net032 net027 net0107 VDD pch_mac l=30n w=100n
MM50_1 ml_b ml_ax VDD VDD pch_mac l=30n w=335.00n
MM50_2 ml_b ml_ax VDD VDD pch_mac l=30n w=335.00n
MM26 net034 D VDD VDD pch_mac l=30n w=170.0n
MM45 ml_ax clkbb net032 VDD pch_mac l=30n w=240.0n
.ENDS
.SUBCKT SDFCNQARD2 SI D SE CP CDN Q VDD VSS
MM3 net89 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM2 qf_x qf net89 VSS nch_mac l=30.0n w=0.14u
MM5 net108 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM7 qf clkb net108 VSS nch_mac l=30.0n w=0.15u
MM52 net109 SE net112 VSS nch_mac l=30.0n w=100n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.15u
MM48 net0220 D VSS VSS nch_mac l=30.0n w=0.175u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net132 mq net133 VSS nch_mac l=30.0n w=100n
MM57 net0219 SE VSS VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net132 VSS nch_mac l=30.0n w=100n
MM66 net133 CDN VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140n
MM46 mq_x clkb net109 VSS nch_mac l=30.0n w=0.165u
MM76 qf_x qf net157 VSS nch_mac l=30.0n w=0.14u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.15u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140n
MM75 net157 CDN VSS VSS nch_mac l=30.0n w=0.14u
MM51 net112 SI VSS VSS nch_mac l=30.0n w=100n
MM47 net109 net0219 net0220 VSS nch_mac l=30.0n w=0.175u
MM1 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u 
MM0 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM0_2 qf_x CDN VDD VDD pch_mac l=30.0n w=0.17u 
MM4 net56 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM42 net25 net0219 net28 VDD pch_mac l=30.0n w=0.12u
MM45 mq_x clkbb net25 VDD pch_mac l=30.0n w=0.22u
MM58 net0219 SE VDD VDD pch_mac l=30.0n w=0.275u
MM60 net76 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net28 SI VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.17u
MM61 net76 mq VDD VDD pch_mac l=30.0n w=120n
MM6 qf clkbb net56 VDD pch_mac l=30.0n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM44 net25 SE net0220 VDD pch_mac l=30.0n w=0.275u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net76 VDD pch_mac l=30.0n w=0.12u
MM43 net0220 D VDD VDD pch_mac l=30.0n w=0.275u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFCNQD2 SI D SE CP CDN Q VDD VSS
MM3 net89 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM2 qf_x qf net89 VSS nch_mac l=30.0n w=245.00n
MM5 net108 qf_x VSS VSS nch_mac l=30.0n w=0.12u
MM7 qf clkb net108 VSS nch_mac l=30.0n w=0.12u
MM52 net109 SE net112 VSS nch_mac l=30.0n w=100n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.155u
MM48 net0220 D VSS VSS nch_mac l=30.0n w=0.175u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net132 mq net133 VSS nch_mac l=30.0n w=100n
MM57 net0219 SE VSS VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net132 VSS nch_mac l=30.0n w=100n
MM66 net133 CDN VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net109 VSS nch_mac l=30.0n w=0.165u
MM76 qf_x qf net157 VSS nch_mac l=30.0n w=0.245u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.245u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM75 net157 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM51 net112 SI VSS VSS nch_mac l=30.0n w=100n
MM47 net109 net0219 net0220 VSS nch_mac l=30.0n w=0.175u
MM1 qf_x qf VDD VDD pch_mac l=30.0n w=0.295u 
MM1_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.295u 
MM0 qf_x CDN VDD VDD pch_mac l=30.0n w=0.12u
MM0B qf_x CDN VDD VDD pch_mac l=30.0n w=0.295u
MM4 net56 qf_x VDD VDD pch_mac l=30.0n w=0.3u
MM42 net25 net0219 net28 VDD pch_mac l=30.0n w=0.12u
MM45 mq_x clkbb net25 VDD pch_mac l=30.0n w=0.22u
MM58 net0219 SE VDD VDD pch_mac l=30.0n w=0.275u
MM60 net76 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net28 SI VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.295u
MM61 net76 mq VDD VDD pch_mac l=30.0n w=120.0n
MM6 qf clkbb net56 VDD pch_mac l=30.0n w=0.12u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM44 net25 SE net0220 VDD pch_mac l=30.0n w=0.275u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net76 VDD pch_mac l=30.0n w=0.12u
MM43 net0220 D VDD VDD pch_mac l=30.0n w=0.275u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFCNQOPTBD2 SI D SE CP CDN Q VDD VSS
MM49_1 ml_b ml_ax VSS VSS nch_mac l=30n w=240.00n
MM49_2 ml_b ml_ax VSS VSS nch_mac l=30n w=240.00n
MM65 net0101 ml_b net0100 VSS nch_mac l=30n w=100n
MM53 clkb CP VSS VSS nch_mac l=30n w=140.0n
MM52 net029 SE net0104 VSS nch_mac l=30n w=100n
MM51 net0104 SI VSS VSS nch_mac l=30n w=100n
MM47_1 net032 D VSS VSS nch_mac l=30n w=135.0n
MM47_2 net032 D VSS VSS nch_mac l=30n w=135.0n
MM64 ml_ax clkbb net0101 VSS nch_mac l=30n w=100n
MM66 net0100 CDN VSS VSS nch_mac l=30n w=100n
MM46 ml_ax clkb net029 VSS nch_mac l=30n w=165.00n
MM55 clkbb clkb VSS VSS nch_mac l=30n w=140.0n
MM75 net0106 CDN VSS VSS nch_mac l=30n w=240.00n
MM76 sl_bx sl_a net0106 VSS nch_mac l=30n w=240.00n
MM71_1 Q sl_bx VSS VSS nch_mac l=30n w=140.0n
MM71_2 Q sl_bx VSS VSS nch_mac l=30n w=140.0n
MM57 net025 SE VSS VSS nch_mac l=30n w=135.0n
MSLTn1 sl_a clkbb ml_b VSS nch_mac l=30n w=155.00n
MM27_1 net029 net025 net032 VSS nch_mac l=30n w=210.0n
MM27_2 net029 net025 net032 VSS nch_mac l=30n w=210.0n
MM7 sl_a clkb net099 VSS nch_mac l=30n w=155.00n
MM5 net099 sl_bx VSS VSS nch_mac l=30n w=140.0n
MM2 sl_bx sl_a net0120 VSS nch_mac l=30n w=240.00n
MM3 net0120 CDN VSS VSS nch_mac l=30n w=240.00n
MM61 net0102 ml_b VDD VDD pch_mac l=30n w=120.0n
MM50_1 ml_b ml_ax VDD VDD pch_mac l=30n w=335.00n
MM50_2 ml_b ml_ax VDD VDD pch_mac l=30n w=335.00n
MM42 net030 net025 net0103 VDD pch_mac l=30n w=100n
MM41 net0103 SI VDD VDD pch_mac l=30n w=100n
MM54 clkb CP VDD VDD pch_mac l=30n w=170.0n
MSLTp1 sl_a clkb ml_b VDD pch_mac l=30n w=295.00n
MM45 ml_ax clkbb net030 VDD pch_mac l=30n w=240.0n
MM72_1 Q sl_bx VDD VDD pch_mac l=30n w=170.0n
MM72_2 Q sl_bx VDD VDD pch_mac l=30n w=170.0n
MM77_1 sl_bx sl_a VDD VDD pch_mac l=30n w=170.0n
MM77_2 sl_bx sl_a VDD VDD pch_mac l=30n w=170.0n
MM78 sl_bx CDN VDD VDD pch_mac l=30n w=170.0n
MM6 sl_a clkbb net0107 VDD pch_mac l=30n w=120.0n
MM56 clkbb clkb VDD VDD pch_mac l=30n w=170.0n
MM17 net032 D VDD VDD pch_mac l=30n w=170.0n
MM4 net0107 sl_bx VDD VDD pch_mac l=30n w=300n
MM26 net032 D VDD VDD pch_mac l=30n w=170.0n
MM60 net0102 CDN VDD VDD pch_mac l=30n w=120.0n
MM58 net025 SE VDD VDD pch_mac l=30n w=170.0n
MM79 ml_ax clkb net0102 VDD pch_mac l=30n w=120.0n
MM44_1 net030 SE net032 VDD pch_mac l=30n w=240.00n
MM44_2 net030 SE net032 VDD pch_mac l=30n w=240.00n
.ENDS
.SUBCKT SDFCSND2 SI D SE CP CDN SDN Q QN VDD VSS
MM6 net0399 SDN net99 VSS nch_mac l=30.0n w=0.155u
MM7 net99 qf_x VSS VSS nch_mac l=30.0n w=0.155u
MM3 net103 SDN VSS VSS nch_mac l=30.0n w=0.22u
MM2 mq mq_x net103 VSS nch_mac l=30.0n w=0.14u
MM52 net111 SE net171 VSS nch_mac l=30.0n w=100n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.155u
MM48 net79 D VSS VSS nch_mac l=30.0n w=0.175u
MM67 net0399 clkb qf VSS nch_mac l=30.0n w=0.155u
MM69 QN net0399 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net0399 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net135 mq net138 VSS nch_mac l=30.0n w=100n
MM57 net0236 SE VSS VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net135 VSS nch_mac l=30.0n w=100n
MM66 net138 CDN VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net111 VSS nch_mac l=30.0n w=0.165u
MM76 qf_x qf net167 VSS nch_mac l=30.0n w=0.22u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM75 net167 CDN VSS VSS nch_mac l=30.0n w=0.22u
MM51 net171 SI VSS VSS nch_mac l=30.0n w=100n
MM47 net111 net0236 net79 VSS nch_mac l=30.0n w=0.175u
MM5 net0399 SDN VDD VDD pch_mac l=30.0n w=0.12u
MM4 net0399 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM42 net19 net0236 net22 VDD pch_mac l=30.0n w=0.12u
MM45 mq_x clkbb net19 VDD pch_mac l=30.0n w=0.22u
MM70 QN net0399 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net0399 VDD VDD pch_mac l=30.0n w=0.17u 
MM58 net0236 SE VDD VDD pch_mac l=30.0n w=0.275u
MM60 net78 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net22 SI VDD VDD pch_mac l=30.0n w=0.12u
MM0 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
MM61 net78 mq VDD VDD pch_mac l=30.0n w=120.0n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM78 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x CDN VDD VDD pch_mac l=30.0n w=0.12u
MM44 net19 SE net79 VDD pch_mac l=30.0n w=0.275u
MM68 net0399 clkbb qf VDD pch_mac l=30.0n w=0.16u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net78 VDD pch_mac l=30.0n w=0.12u
MM43 net79 D VDD VDD pch_mac l=30.0n w=0.275u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM1 mq mq_x VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFCSNQD2 SI D SE CP CDN SDN Q VDD VSS
MM10 net0109 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM11 qf_x qf net0109 VSS nch_mac l=30.0n w=0.245u
MM47 net86 net0245 net130 VSS nch_mac l=30.0n w=0.175u
MM51 net89 SI VSS VSS nch_mac l=30.0n w=100n
MM75 net49 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM76 qf_x qf net49 VSS nch_mac l=30.0n w=0.245u
MM46 mq_x clkb net86 VSS nch_mac l=30.0n w=0.165u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM66 net58 CDN VSS VSS nch_mac l=30.0n w=100n
MM64 mq_x clkbb net65 VSS nch_mac l=30.0n w=100n
MM57 net0245 SE VSS VSS nch_mac l=30.0n w=0.12u
MM65 net65 mq net58 VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net0163 clkb qf VSS nch_mac l=30.0n w=0.155u
MM48 net130 D VSS VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.155u
MM52 net86 SE net89 VSS nch_mac l=30.0n w=100n
MM2 mq mq_x net94 VSS nch_mac l=30.0n w=0.14u
MM3 net94 SDN VSS VSS nch_mac l=30.0n w=0.245u
MM7 net29 qf_x VSS VSS nch_mac l=30.0n w=0.155u
MM6 net0163 SDN net29 VSS nch_mac l=30.0n w=0.155u
MM8 qf_x CDN VDD VDD pch_mac l=30.0n w=0.12u
MM8B qf_x CDN VDD VDD pch_mac l=30.0n w=0.315u
MM1 mq mq_x VDD VDD pch_mac l=30.0n w=0.17u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM43 net130 D VDD VDD pch_mac l=30.0n w=0.275u
MM79 mq_x clkb net137 VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net0163 clkbb qf VDD pch_mac l=30.0n w=0.16u
MM44 net182 SE net130 VDD pch_mac l=30.0n w=0.275u
MM78 qf_x qf VDD VDD pch_mac l=30.0n w=0.315u 
MM78_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.315u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM61 net137 mq VDD VDD pch_mac l=30.0n w=120.0n
MM0 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net166 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net137 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM58 net0245 SE VDD VDD pch_mac l=30.0n w=0.275u
MM45 mq_x clkbb net182 VDD pch_mac l=30.0n w=0.22u
MM42 net182 net0245 net166 VDD pch_mac l=30.0n w=0.12u
MM4 net0163 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM5 net0163 SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFD2 SI D SE CP Q QN VDD VSS
MM73 net101 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM69 QN net101 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net101 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 qf_x qf VSS VSS nch_mac l=30.0n w=0.14u
MM52 net89 SE net92 VSS nch_mac l=30.0n w=100n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.265u
MM48 net0268 D VSS VSS nch_mac l=30.0n w=0.175u
MM67 net101 clkb qf VSS nch_mac l=30.0n w=0.265u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 mq_x clkbb net112 VSS nch_mac l=30.0n w=100n
MM57 net0196 SE VSS VSS nch_mac l=30.0n w=0.175u
MM66 net112 mq VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net89 VSS nch_mac l=30.0n w=0.175u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.265u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM51 net92 SI VSS VSS nch_mac l=30.0n w=100n
MM47 net89 net0196 net0268 VSS nch_mac l=30.0n w=0.175u
MM70 QN net101 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net101 VDD VDD pch_mac l=30.0n w=0.17u 
MM74 net101 qf_x VDD VDD pch_mac l=30.0n w=0.335u
MM1 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u
MM0 mq_x clkb net0107 VDD pch_mac l=30.0n w=0.12u
MM42 net25 net0196 net37 VDD pch_mac l=30.0n w=0.12u
MM45 mq_x clkbb net25 VDD pch_mac l=30.0n w=200n
MM58 net0196 SE VDD VDD pch_mac l=30.0n w=0.24u
MM41 net37 SI VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.285u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM44 net25 SE net0268 VDD pch_mac l=30.0n w=0.24u
MM68 net101 clkbb qf VDD pch_mac l=30.0n w=0.285u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 net0107 mq VDD VDD pch_mac l=30.0n w=100n
MM43 net0268 D VDD VDD pch_mac l=30.0n w=0.24u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.285u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFKCNARD2 SI D SE CP CN Q QN VDD VSS
MM13 net86 SI VSS VSS nch_mac l=30.0n w=0.145u
MM16 net90 SE VSS VSS nch_mac l=30.0n w=0.145u
MM1 net94 CN net98 VSS nch_mac l=30.0n w=0.145u
MM3 net98 D VSS VSS nch_mac l=30.0n w=0.14u
MM6 net42 net90 net94 VSS nch_mac l=30.0n w=0.145u
MM12 net42 SE net86 VSS nch_mac l=30.0n w=0.145u
MM20 mq clkb net30 VSS nch_mac l=30.0n w=0.15u
MM9 net121 qf VSS VSS nch_mac l=30.0n w=0.15u
MM10 qf_x clkb net121 VSS nch_mac l=30.0n w=0.15u
MM18 net30 net42 VSS VSS nch_mac l=30.0n w=0.15u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.15u
MM69 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net149 mq_x VSS VSS nch_mac l=30.0n w=0.15u
MM64 mq clkbb net149 VSS nch_mac l=30.0n w=0.15u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.15u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140n
MM14 net45 SI VDD VDD pch_mac l=30.0n w=0.185u
MM5 net42 SE net94 VDD pch_mac l=30.0n w=0.185u
MM15 net90 SE VDD VDD pch_mac l=30.0n w=0.17u
MM7 net22 qf VDD VDD pch_mac l=30.0n w=0.17u
MM19 mq clkbb net30 VDD pch_mac l=30.0n w=0.215u
MM17 net30 net42 VDD VDD pch_mac l=30.0n w=0.215u
MM4 net94 CN VDD VDD pch_mac l=30.0n w=0.185u
MM8 qf_x clkbb net22 VDD pch_mac l=30.0n w=0.17u
MM11 net42 net90 net45 VDD pch_mac l=30.0n w=0.185u
MM2 net94 D VDD VDD pch_mac l=30.0n w=0.17u
MM70 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net58 mq_x VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq clkb net58 VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.17u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFKCND2 SI D SE CP CN Q QN VDD VSS
MM13 net86 SI VSS VSS nch_mac l=30.0n w=0.145u
MM16 net90 SE VSS VSS nch_mac l=30.0n w=0.145u
MM1 net94 CN net98 VSS nch_mac l=30.0n w=0.145u
MM3 net98 D VSS VSS nch_mac l=30.0n w=0.14u
MM6 net42 net90 net94 VSS nch_mac l=30.0n w=0.145u
MM12 net42 SE net86 VSS nch_mac l=30.0n w=0.145u
MM20 mq clkb net30 VSS nch_mac l=30.0n w=0.155u
MM9 net121 qf VSS VSS nch_mac l=30.0n w=0.12u
MM10 qf_x clkb net121 VSS nch_mac l=30.0n w=0.12u
MM18 net30 net42 VSS VSS nch_mac l=30.0n w=0.155u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.265u
MM69 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net149 mq_x VSS VSS nch_mac l=30.0n w=100n
MM64 mq clkbb net149 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.18u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM14 net45 SI VDD VDD pch_mac l=30.0n w=0.185u
MM5 net42 SE net94 VDD pch_mac l=30.0n w=0.185u
MM15 net90 SE VDD VDD pch_mac l=30.0n w=0.17u
MM7 net22 qf VDD VDD pch_mac l=30.0n w=0.12u
MM19 mq clkbb net30 VDD pch_mac l=30.0n w=0.215u
MM17 net30 net42 VDD VDD pch_mac l=30.0n w=0.215u
MM4 net94 CN VDD VDD pch_mac l=30.0n w=0.185u
MM8 qf_x clkbb net22 VDD pch_mac l=30.0n w=0.275u
MM11 net42 net90 net45 VDD pch_mac l=30.0n w=0.185u
MM2 net94 D VDD VDD pch_mac l=30.0n w=0.17u
MM70 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net58 mq_x VDD VDD pch_mac l=30.0n w=100n
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq clkb net58 VDD pch_mac l=30.0n w=100n
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFKCNQARD2 SI D SE CP CN Q VDD VSS
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.15u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140n
MM64 mq clkbb net25 VSS nch_mac l=30.0n w=0.15u
MM65 net25 mq_x VSS VSS nch_mac l=30.0n w=0.15u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.15u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM18 net129 net57 VSS VSS nch_mac l=30.0n w=0.15u
MM10 qf_x clkb net49 VSS nch_mac l=30.0n w=0.15u
MM9 net49 qf VSS VSS nch_mac l=30.0n w=0.15u
MM20 mq clkb net129 VSS nch_mac l=30.0n w=0.15u
MM12 net57 SE net77 VSS nch_mac l=30.0n w=0.145u
MM6 net57 net141 net69 VSS nch_mac l=30.0n w=0.145u
MM3 net65 D VSS VSS nch_mac l=30.0n w=0.14u
MM1 net69 CN net65 VSS nch_mac l=30.0n w=0.145u
MM16 net141 SE VSS VSS nch_mac l=30.0n w=0.145u
MM13 net77 SI VSS VSS nch_mac l=30.0n w=0.145u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.185u
MM79 mq clkb net92 VDD pch_mac l=30.0n w=0.185u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.185u
MM60 net92 mq_x VDD VDD pch_mac l=30.0n w=0.185u
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM2 net69 D VDD VDD pch_mac l=30.0n w=0.17u
MM11 net57 net141 net120 VDD pch_mac l=30.0n w=0.185u
MM8 qf_x clkbb net137 VDD pch_mac l=30.0n w=0.185u
MM4 net69 CN VDD VDD pch_mac l=30.0n w=0.185u
MM17 net129 net57 VDD VDD pch_mac l=30.0n w=0.215u
MM19 mq clkbb net129 VDD pch_mac l=30.0n w=0.215u
MM7 net137 qf VDD VDD pch_mac l=30.0n w=0.185u
MM15 net141 SE VDD VDD pch_mac l=30.0n w=0.17u
MM5 net57 SE net69 VDD pch_mac l=30.0n w=0.185u
MM14 net120 SI VDD VDD pch_mac l=30.0n w=0.185u
.ENDS
.SUBCKT SDFKCNQD2 SI D SE CP CN Q VDD VSS
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.18u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM64 mq clkbb net25 VSS nch_mac l=30.0n w=100n
MM65 net25 mq_x VSS VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.265u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM18 net129 net57 VSS VSS nch_mac l=30.0n w=0.155u
MM10 qf_x clkb net49 VSS nch_mac l=30.0n w=0.12u
MM9 net49 qf VSS VSS nch_mac l=30.0n w=0.12u
MM20 mq clkb net129 VSS nch_mac l=30.0n w=0.155u
MM12 net57 SE net77 VSS nch_mac l=30.0n w=0.145u
MM6 net57 net141 net69 VSS nch_mac l=30.0n w=0.145u
MM3 net65 D VSS VSS nch_mac l=30.0n w=0.14u
MM1 net69 CN net65 VSS nch_mac l=30.0n w=0.145u
MM16 net141 SE VSS VSS nch_mac l=30.0n w=0.145u
MM13 net77 SI VSS VSS nch_mac l=30.0n w=0.145u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.275u
MM79 mq clkb net92 VDD pch_mac l=30.0n w=100n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.275u
MM60 net92 mq_x VDD VDD pch_mac l=30.0n w=100n
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM2 net69 D VDD VDD pch_mac l=30.0n w=0.17u
MM11 net57 net141 net120 VDD pch_mac l=30.0n w=0.185u
MM8 qf_x clkbb net137 VDD pch_mac l=30.0n w=0.275u
MM4 net69 CN VDD VDD pch_mac l=30.0n w=0.185u
MM17 net129 net57 VDD VDD pch_mac l=30.0n w=0.215u
MM19 mq clkbb net129 VDD pch_mac l=30.0n w=0.215u
MM7 net137 qf VDD VDD pch_mac l=30.0n w=0.12u
MM15 net141 SE VDD VDD pch_mac l=30.0n w=0.17u
MM5 net57 SE net69 VDD pch_mac l=30.0n w=0.185u
MM14 net120 SI VDD VDD pch_mac l=30.0n w=0.185u
.ENDS
.SUBCKT SDFKCSND2 SI D SE CP CN SN Q QN VDD VSS
MM22 net99 SN VSS VSS nch_mac l=30.0n w=0.245u
MM0 net83 net99 net86 VSS nch_mac l=30.0n w=0.12u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.18u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM64 mq clkbb net35 VSS nch_mac l=30.0n w=100n
MM65 net35 mq_x VSS VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM69 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.265u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM18 net155 net143 VSS VSS nch_mac l=30.0n w=0.155u
MM10 qf_x clkb net63 VSS nch_mac l=30.0n w=0.12u
MM9 net63 qf VSS VSS nch_mac l=30.0n w=0.12u
MM20 mq clkb net155 VSS nch_mac l=30.0n w=0.155u
MM12 net143 SE net91 VSS nch_mac l=30.0n w=0.12u
MM6 net143 net87 net83 VSS nch_mac l=30.0n w=0.215u
MM3 net86 CN VSS VSS nch_mac l=30.0n w=0.245u
MM1 net83 D net86 VSS nch_mac l=30.0n w=0.245u
MM16 net87 SE VSS VSS nch_mac l=30.0n w=0.12u
MM13 net91 SI VSS VSS nch_mac l=30.0n w=0.12u
MM21 net142 net99 VDD VDD pch_mac l=30.0n w=0.205u
MM23 net99 SN VDD VDD pch_mac l=30.0n w=0.12u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.275u
MM79 mq clkb net114 VDD pch_mac l=30.0n w=100n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.275u
MM60 net114 mq_x VDD VDD pch_mac l=30.0n w=100n
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM70 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM2 net83 D net142 VDD pch_mac l=30.0n w=0.205u
MM11 net143 net87 net146 VDD pch_mac l=30.0n w=0.12u
MM8 qf_x clkbb net163 VDD pch_mac l=30.0n w=0.275u
MM4 net83 CN VDD VDD pch_mac l=30.0n w=0.12u
MM17 net155 net143 VDD VDD pch_mac l=30.0n w=0.215u
MM19 mq clkbb net155 VDD pch_mac l=30.0n w=0.215u
MM7 net163 qf VDD VDD pch_mac l=30.0n w=0.12u
MM15 net87 SE VDD VDD pch_mac l=30.0n w=0.17u
MM5 net143 SE net83 VDD pch_mac l=30.0n w=0.195u
MM14 net146 SI VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFKCSNQD2 SI D SE CP CN SN Q VDD VSS
MM13 net113 SI VSS VSS nch_mac l=30.0n w=0.12u
MM16 net201 SE VSS VSS nch_mac l=30.0n w=0.12u
MM1 net121 D net125 VSS nch_mac l=30.0n w=0.245u
MM3 net125 CN VSS VSS nch_mac l=30.0n w=0.245u
MM6 net225 net201 net121 VSS nch_mac l=30.0n w=0.215u
MM12 net225 SE net113 VSS nch_mac l=30.0n w=0.12u
MM20 mq clkb net213 VSS nch_mac l=30.0n w=0.155u
MM9 net148 qf VSS VSS nch_mac l=30.0n w=0.12u
MM10 qf_x clkb net148 VSS nch_mac l=30.0n w=0.12u
MM18 net213 net225 VSS VSS nch_mac l=30.0n w=0.155u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.265u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net165 mq_x VSS VSS nch_mac l=30.0n w=100n
MM64 mq clkbb net165 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.18u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM0 net121 net265 net125 VSS nch_mac l=30.0n w=0.12u
MM22 net265 SN VSS VSS nch_mac l=30.0n w=0.245u
MM14 net228 SI VDD VDD pch_mac l=30.0n w=0.12u
MM5 net225 SE net121 VDD pch_mac l=30.0n w=0.195u
MM15 net201 SE VDD VDD pch_mac l=30.0n w=0.17u
MM7 net224 qf VDD VDD pch_mac l=30.0n w=0.12u
MM19 mq clkbb net213 VDD pch_mac l=30.0n w=0.215u
MM17 net213 net225 VDD VDD pch_mac l=30.0n w=0.215u
MM4 net121 CN VDD VDD pch_mac l=30.0n w=0.12u
MM8 qf_x clkbb net224 VDD pch_mac l=30.0n w=0.275u
MM11 net225 net201 net228 VDD pch_mac l=30.0n w=0.12u
MM2 net121 D net232 VDD pch_mac l=30.0n w=0.205u
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net256 mq_x VDD VDD pch_mac l=30.0n w=100n
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq clkb net256 VDD pch_mac l=30.0n w=100n
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM23 net265 SN VDD VDD pch_mac l=30.0n w=0.12u
MM21 net232 net265 VDD VDD pch_mac l=30.0n w=0.205u
.ENDS
.SUBCKT SDFKSND2 SI D SE CP SN Q QN VDD VSS
MM13 net90 SI VSS VSS nch_mac l=30.0n w=0.12u
MM16 net94 SE VSS VSS nch_mac l=30.0n w=0.12u
MM1 net98 D VSS VSS nch_mac l=30.0n w=0.14u
MM6 net38 net94 net98 VSS nch_mac l=30.0n w=0.26u
MM12 net38 SE net90 VSS nch_mac l=30.0n w=0.12u
MM20 mq clkb net30 VSS nch_mac l=30.0n w=0.155u
MM9 net114 qf VSS VSS nch_mac l=30.0n w=0.12u
MM10 qf_x clkb net114 VSS nch_mac l=30.0n w=0.12u
MM18 net30 net38 VSS VSS nch_mac l=30.0n w=0.155u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.265u
MM69 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net149 mq_x VSS VSS nch_mac l=30.0n w=100n
MM64 mq clkbb net149 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.18u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM0 net98 net166 VSS VSS nch_mac l=30.0n w=0.14u
MM22 net166 SN VSS VSS nch_mac l=30.0n w=0.14u
MM14 net10 SI VDD VDD pch_mac l=30.0n w=0.12u
MM5 net38 SE net98 VDD pch_mac l=30.0n w=0.3u
MM15 net94 SE VDD VDD pch_mac l=30.0n w=0.17u
MM7 net37 qf VDD VDD pch_mac l=30.0n w=0.12u
MM19 mq clkbb net30 VDD pch_mac l=30.0n w=0.215u
MM17 net30 net38 VDD VDD pch_mac l=30.0n w=0.215u
MM8 qf_x clkbb net37 VDD pch_mac l=30.0n w=0.275u
MM11 net38 net94 net10 VDD pch_mac l=30.0n w=0.12u
MM2 net98 D net86 VDD pch_mac l=30.0n w=0.3u
MM70 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM60 net73 mq_x VDD VDD pch_mac l=30.0n w=100n
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq clkb net73 VDD pch_mac l=30.0n w=100n
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.275u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM23 net166 SN VDD VDD pch_mac l=30.0n w=0.12u
MM21 net86 net166 VDD VDD pch_mac l=30.0n w=0.3u
.ENDS
.SUBCKT SDFKSNQD2 SI D SE CP SN Q VDD VSS
MM22 net9 SN VSS VSS nch_mac l=30.0n w=0.14u
MM0 net73 net9 VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.18u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM64 mq clkbb net33 VSS nch_mac l=30.0n w=100n
MM65 net33 mq_x VSS VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.265u
MM73 qf qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM18 net49 net65 VSS VSS nch_mac l=30.0n w=0.155u
MM10 qf_x clkb net57 VSS nch_mac l=30.0n w=0.12u
MM9 net57 qf VSS VSS nch_mac l=30.0n w=0.12u
MM20 mq clkb net49 VSS nch_mac l=30.0n w=0.155u
MM12 net65 SE net68 VSS nch_mac l=30.0n w=0.12u
MM6 net65 net77 net73 VSS nch_mac l=30.0n w=0.26u
MM1 net73 D VSS VSS nch_mac l=30.0n w=0.14u
MM16 net77 SE VSS VSS nch_mac l=30.0n w=0.12u
MM13 net68 SI VSS VSS nch_mac l=30.0n w=0.12u
MM21 net85 net9 VDD VDD pch_mac l=30.0n w=0.3u
MM23 net9 SN VDD VDD pch_mac l=30.0n w=0.12u
MM54 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.275u
MM79 mq clkb net104 VDD pch_mac l=30.0n w=100n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.275u
MM60 net104 mq_x VDD VDD pch_mac l=30.0n w=100n
MM74 qf qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM2 net73 D net85 VDD pch_mac l=30.0n w=0.3u
MM11 net65 net77 net157 VDD pch_mac l=30.0n w=0.12u
MM8 qf_x clkbb net136 VDD pch_mac l=30.0n w=0.275u
MM17 net49 net65 VDD VDD pch_mac l=30.0n w=0.215u
MM19 mq clkbb net49 VDD pch_mac l=30.0n w=0.215u
MM7 net136 qf VDD VDD pch_mac l=30.0n w=0.12u
MM15 net77 SE VDD VDD pch_mac l=30.0n w=0.17u
MM5 net65 SE net73 VDD pch_mac l=30.0n w=0.3u
MM14 net157 SI VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFMD2 DA DB SA SI SE CP Q QN VDD VSS
MSLTn1 qf_x clkbb net0413 VSS nch_mac l=30.0n w=0.14u
MSLTn2 net0413 mq VSS VSS nch_mac l=30.0n w=0.14u
MM16 net0402 qf VSS VSS nch_mac l=30.0n w=0.12u
MM47 net167 DA net102 VSS nch_mac l=30.0n w=0.22u
MM51 net103 SI VSS VSS nch_mac l=30.0n w=100n
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.275u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.195u
MM76 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net167 VSS nch_mac l=30.0n w=0.27u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.195u
MM64 mq_x clkbb net139 VSS nch_mac l=30.0n w=100n
MM57 net63 SE VSS VSS nch_mac l=30.0n w=0.12u
MM65 net139 mq VSS VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM15 qf_x clkb net0402 VSS nch_mac l=30.0n w=0.12u
MM48 net102 SA net182 VSS nch_mac l=30.0n w=0.22u
MM73 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM73_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM52 net167 SE net103 VSS nch_mac l=30.0n w=100n
MM7 net182 net63 VSS VSS nch_mac l=30.0n w=0.185u
MM0 net175 SA VSS VSS nch_mac l=30.0n w=0.14u
MM3 net179 DB net182 VSS nch_mac l=30.0n w=0.185u
MM2 net167 net175 net179 VSS nch_mac l=30.0n w=0.22u
MM13 qf_x clkbb net0325 VDD pch_mac l=30.0n w=0.12u
MSLTp1 net0330 mq VDD VDD pch_mac l=30.0n w=0.31u
MSLTp2 qf_x clkb net0330 VDD pch_mac l=30.0n w=0.31u
MM43 net15 net175 net86 VDD pch_mac l=30.0n w=0.175u
MM79 mq_x clkb net55 VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM14 net0325 qf VDD VDD pch_mac l=30.0n w=0.12u
MM44 net79 DA net15 VDD pch_mac l=30.0n w=0.175u
MM77 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=170.0n
MM41 net51 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net55 mq VDD VDD pch_mac l=30.0n w=0.12u
MM74 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM74_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM58 net63 SE VDD VDD pch_mac l=30.0n w=0.14u
MM45 mq_x clkbb net79 VDD pch_mac l=30.0n w=0.21u
MM6 net86 SE VDD VDD pch_mac l=30.0n w=0.22u
MM42 net79 net63 net51 VDD pch_mac l=30.0n w=0.12u
MM5 net90 DB net86 VDD pch_mac l=30.0n w=0.22u
MM4 net79 SA net90 VDD pch_mac l=30.0n w=0.175u
MM1 net175 SA VDD VDD pch_mac l=30.0n w=0.17u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.305u
.ENDS
.SUBCKT SDFMQD2 DA DB SA SI SE CP Q VDD VSS
MM2 net26 net98 net14 VSS nch_mac l=30.0n w=0.22u
MM3 net14 DB net17 VSS nch_mac l=30.0n w=0.185u
MM0 net98 SA VSS VSS nch_mac l=30.0n w=0.14u
MM7 net17 net122 VSS VSS nch_mac l=30.0n w=0.185u
MM52 net26 SE net74 VSS nch_mac l=30.0n w=100n
MM48 net81 SA net17 VSS nch_mac l=30.0n w=0.22u
MM15 qf_x clkb net82 VSS nch_mac l=30.0n w=0.12u
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net42 mq VSS VSS nch_mac l=30.0n w=100n
MM57 net122 SE VSS VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkbb net42 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.195u
MM46 mq_x clkb net26 VSS nch_mac l=30.0n w=0.27u
MM76 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.195u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.275u
MM51 net74 SI VSS VSS nch_mac l=30.0n w=100n
MM47 net26 DA net81 VSS nch_mac l=30.0n w=0.22u
MM16 net82 qf VSS VSS nch_mac l=30.0n w=0.12u
MSLTn2 net93 mq VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf_x clkbb net93 VSS nch_mac l=30.0n w=0.14u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.305u
MM1 net98 SA VDD VDD pch_mac l=30.0n w=0.17u
MM4 net110 SA net120 VDD pch_mac l=30.0n w=0.175u
MM5 net120 DB net109 VDD pch_mac l=30.0n w=0.22u
MM42 net110 net122 net130 VDD pch_mac l=30.0n w=0.12u
MM6 net109 SE VDD VDD pch_mac l=30.0n w=0.22u
MM45 mq_x clkbb net110 VDD pch_mac l=30.0n w=0.21u
MM58 net122 SE VDD VDD pch_mac l=30.0n w=0.14u
MM60 net161 mq VDD VDD pch_mac l=30.0n w=0.12u
MM41 net130 SI VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=170.0n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM44 net110 DA net149 VDD pch_mac l=30.0n w=0.175u
MM14 net177 qf VDD VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net161 VDD pch_mac l=30.0n w=0.12u
MM43 net149 net98 net109 VDD pch_mac l=30.0n w=0.175u
MSLTp2 qf_x clkb net170 VDD pch_mac l=30.0n w=0.31u
MSLTp1 net170 mq VDD VDD pch_mac l=30.0n w=0.31u
MM13 qf_x clkbb net177 VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFNCND2 SI D SE CPN CDN Q QN VDD VSS
MM5 net0188 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM4 qf_x qf net0188 VSS nch_mac l=30.0n w=0.245u
MM52 net86 SE net89 VSS nch_mac l=30.0n w=100n
MM73 net102 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.155u
MM48 net74 D VSS VSS nch_mac l=30.0n w=0.175u
MM67 net102 clkbb qf VSS nch_mac l=30.0n w=0.155u
MM69 QN net102 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net102 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net125 mq net117 VSS nch_mac l=30.0n w=100n
MM57 net0209 SE VSS VSS nch_mac l=30.0n w=0.12u
MM64 mq_x clkb net125 VSS nch_mac l=30.0n w=100n
MM66 net117 CDN VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkbb net86 VSS nch_mac l=30.0n w=0.165u
MM76 qf_x qf net141 VSS nch_mac l=30.0n w=0.245u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.245u
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=140.0n
MM75 net141 CDN VSS VSS nch_mac l=30.0n w=0.245u
MM47 net86 net0209 net74 VSS nch_mac l=30.0n w=0.175u
MM80 net89 SI VSS VSS nch_mac l=30.0n w=0.12u
MM0 qf_x CDN VDD VDD pch_mac l=30.0n w=0.12u
MM0B qf_x CDN VDD VDD pch_mac l=30.0n w=0.295u
MM42 net10 net0209 net34 VDD pch_mac l=30.0n w=0.12u
MM45 mq_x clkb net10 VDD pch_mac l=30.0n w=0.22u
MM70 QN net102 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net102 VDD VDD pch_mac l=30.0n w=0.17u 
MM58 net0209 SE VDD VDD pch_mac l=30.0n w=0.275u
MM74 net102 qf_x VDD VDD pch_mac l=30.0n w=0.3u
MM60 net30 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net34 SI VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.295u
MM61 net30 mq VDD VDD pch_mac l=30.0n w=120.0n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=0.295u 
MM77_2 qf_x qf VDD VDD pch_mac l=30.0n w=0.295u 
MM44 net10 SE net74 VDD pch_mac l=30.0n w=0.275u
MM68 net102 clkb qf VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkbb net30 VDD pch_mac l=30.0n w=0.12u
MM43 net74 D VDD VDD pch_mac l=30.0n w=0.275u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.295u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFNCSND2 SI D SE CPN CDN SDN Q QN VDD VSS
MM47 net75 net0253 net67 VSS nch_mac l=30.0n w=0.175u
MM51 net78 SI VSS VSS nch_mac l=30.0n w=100n
MM75 net30 CDN VSS VSS nch_mac l=30.0n w=0.22u
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=140.0n
MM76 qf_x qf net30 VSS nch_mac l=30.0n w=0.22u
MM46 mq_x clkbb net75 VSS nch_mac l=30.0n w=0.165u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM66 net54 CDN VSS VSS nch_mac l=30.0n w=100n
MM64 mq_x clkb net51 VSS nch_mac l=30.0n w=100n
MM57 net0253 SE VSS VSS nch_mac l=30.0n w=0.12u
MM65 net51 mq net54 VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM69 QN net0161 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net0161 VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net0161 clkbb qf VSS nch_mac l=30.0n w=0.155u
MM48 net67 D VSS VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.155u
MM52 net75 SE net78 VSS nch_mac l=30.0n w=100n
MM2 mq mq_x net83 VSS nch_mac l=30.0n w=0.14u
MM3 net83 SDN VSS VSS nch_mac l=30.0n w=0.22u
MM7 net94 qf_x VSS VSS nch_mac l=30.0n w=0.155u
MM6 net0161 SDN net94 VSS nch_mac l=30.0n w=0.155u
MM1 mq mq_x VDD VDD pch_mac l=30.0n w=0.17u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.275u
MM43 net67 D VDD VDD pch_mac l=30.0n w=0.275u
MM79 mq_x clkbb net151 VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net0161 clkb qf VDD pch_mac l=30.0n w=0.16u
MM44 net167 SE net67 VDD pch_mac l=30.0n w=0.275u
MM77 qf_x CDN VDD VDD pch_mac l=30.0n w=0.12u
MM78 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM61 net151 mq VDD VDD pch_mac l=30.0n w=120.0n
MM0 mq SDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net170 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net151 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM58 net0253 SE VDD VDD pch_mac l=30.0n w=0.275u
MM70 QN net0161 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net0161 VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkb net167 VDD pch_mac l=30.0n w=0.22u
MM42 net167 net0253 net170 VDD pch_mac l=30.0n w=0.12u
MM4 net0161 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM5 net0161 SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFND2 SI D SE CPN Q QN VDD VSS
MM47 net69 net0208 net108 VSS nch_mac l=30.0n w=0.175u
MM51 net72 SI VSS VSS nch_mac l=30.0n w=100n
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.265u
MM46 mq_x clkbb net69 VSS nch_mac l=30.0n w=0.175u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM66 net44 mq VSS VSS nch_mac l=30.0n w=100n
MM57 net0208 SE VSS VSS nch_mac l=30.0n w=0.175u
MM65 mq_x clkb net44 VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM69 QN net53 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net53 VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net53 clkbb qf VSS nch_mac l=30.0n w=0.265u
MM48 net108 D VSS VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.265u
MM73 net53 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM52 net69 SE net72 VSS nch_mac l=30.0n w=100n
MM2 qf_x qf VSS VSS nch_mac l=30.0n w=0.14u
MM0 mq_x clkbb net0163 VDD pch_mac l=30.0n w=0.12u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.285u
MM43 net108 D VDD VDD pch_mac l=30.0n w=0.24u
MM79 net0163 mq VDD VDD pch_mac l=30.0n w=100n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net53 clkb qf VDD pch_mac l=30.0n w=0.285u
MM44 net137 SE net108 VDD pch_mac l=30.0n w=0.24u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.285u
MM41 net140 SI VDD VDD pch_mac l=30.0n w=0.12u
MM74 net53 qf_x VDD VDD pch_mac l=30.0n w=0.335u
MM58 net0208 SE VDD VDD pch_mac l=30.0n w=0.24u
MM70 QN net53 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net53 VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkb net137 VDD pch_mac l=30.0n w=200n
MM42 net137 net0208 net140 VDD pch_mac l=30.0n w=0.12u
MM1 qf_x qf VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SDFNSND2 SI D SE CPN SDN Q QN VDD VSS
MM47 net165 net237 net0227 VSS nch_mac l=30.0n w=0.175u
MM51 net113 SI VSS VSS nch_mac l=30.0n w=100n
MM53 clkb CPN VSS VSS nch_mac l=30.0n w=140.0n
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkbb net165 VSS nch_mac l=30.0n w=0.175u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM64 mq_x clkb net136 VSS nch_mac l=30.0n w=100n
MM57 net237 SE VSS VSS nch_mac l=30.0n w=0.12u
MM65 net136 mq VSS VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM69 QN net153 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net153 VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net153 clkbb qf VSS nch_mac l=30.0n w=0.22u
MM48 net0227 D VSS VSS nch_mac l=30.0n w=0.175u
MSLTn1 qf clkb mq VSS nch_mac l=30.0n w=0.22u
MM52 net165 SE net113 VSS nch_mac l=30.0n w=100n
MM2 mq SDN net173 VSS nch_mac l=30.0n w=0.22u
MM3 net173 mq_x VSS VSS nch_mac l=30.0n w=0.22u
MM7 net184 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM6 net153 SDN net184 VSS nch_mac l=30.0n w=0.14u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM1 mq SDN VDD VDD pch_mac l=30.0n w=0.215u
MM54 clkb CPN VDD VDD pch_mac l=30.0n w=0.17u
MSLTp1 qf clkbb mq VDD pch_mac l=30.0n w=0.31u
MM43 net0227 D VDD VDD pch_mac l=30.0n w=0.275u
MM79 mq_x clkbb net208 VDD pch_mac l=30.0n w=100n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net153 clkb qf VDD pch_mac l=30.0n w=0.12u
MM44 net249 SE net0227 VDD pch_mac l=30.0n w=0.275u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM0 mq mq_x VDD VDD pch_mac l=30.0n w=0.215u
MM41 net252 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net208 mq VDD VDD pch_mac l=30.0n w=100n
MM58 net237 SE VDD VDD pch_mac l=30.0n w=0.275u
MM70 QN net153 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net153 VDD VDD pch_mac l=30.0n w=0.17u 
MM45 mq_x clkb net249 VDD pch_mac l=30.0n w=0.22u
MM42 net249 net237 net252 VDD pch_mac l=30.0n w=0.12u
MM4 net153 qf_x VDD VDD pch_mac l=30.0n w=0.17u
MM5 net153 SDN VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFOPTBD2 SI D SE CP Q QN VDD VSS
MM65 ml_ax clkbb net092 VSS nch_mac l=30n w=100n
MM66 net092 ml_b VSS VSS nch_mac l=30n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30n w=140.0n
MM53 clkb CP VSS VSS nch_mac l=30n w=140.0n
MM52 net027 SE net095 VSS nch_mac l=30n w=100n
MM57 net023 SE VSS VSS nch_mac l=30n w=135.0n
MM47_1 net030 D VSS VSS nch_mac l=30n w=135.0n
MM47_2 net030 D VSS VSS nch_mac l=30n w=135.0n
MM51 net095 SI VSS VSS nch_mac l=30n w=100n
MM27_1 net027 net023 net030 VSS nch_mac l=30n w=210.0n
MM27_2 net027 net023 net030 VSS nch_mac l=30n w=210.0n
MM46 ml_ax clkb net027 VSS nch_mac l=30n w=200n
MM15 ml_b ml_ax VSS VSS nch_mac l=30n w=140.0n
MM71_1 Q sl_bx VSS VSS nch_mac l=30n w=140.0n
MM71_2 Q sl_bx VSS VSS nch_mac l=30n w=140.0n
MM67 net101 clkb sl_a VSS nch_mac l=30n w=265.00n
MSLTn1 sl_a clkbb ml_b VSS nch_mac l=30n w=265.00n
MM49 ml_b ml_ax VSS VSS nch_mac l=30n w=140.0n
MM2 sl_bx sl_a VSS VSS nch_mac l=30n w=140.0n
MM69_1 QN net101 VSS VSS nch_mac l=30n w=140.0n
MM69_2 QN net101 VSS VSS nch_mac l=30n w=140.0n
MM73 net101 sl_bx VSS VSS nch_mac l=30n w=140.0n
MM0 ml_ax clkb net093 VDD pch_mac l=30n w=100n
MM79 net093 ml_b VDD VDD pch_mac l=30n w=100n
MM56 clkbb clkb VDD VDD pch_mac l=30n w=325.00n
MM54 clkb CP VDD VDD pch_mac l=30n w=170.0n
MSLTp1 sl_a clkb ml_b VDD pch_mac l=30n w=285.00n
MM58 net023 SE VDD VDD pch_mac l=30n w=170.0n
MM72_1 Q sl_bx VDD VDD pch_mac l=30n w=170.0n
MM72_2 Q sl_bx VDD VDD pch_mac l=30n w=170.0n
MM68 net101 clkbb sl_a VDD pch_mac l=30n w=285.00n
MM50_1 ml_b ml_ax VDD VDD pch_mac l=30n w=325.00n
MM50_2 ml_b ml_ax VDD VDD pch_mac l=30n w=325.00n
MM45 ml_ax clkbb net028 VDD pch_mac l=30n w=200n
MM26 net030 D VDD VDD pch_mac l=30n w=170.0n
MM1 sl_bx sl_a VDD VDD pch_mac l=30n w=170.0n
MM74 net101 sl_bx VDD VDD pch_mac l=30n w=330.0n
MM70_1 QN net101 VDD VDD pch_mac l=30n w=170.0n
MM70_2 QN net101 VDD VDD pch_mac l=30n w=170.0n
MM17 net030 D VDD VDD pch_mac l=30n w=170.0n
MM42 net028 net023 net094 VDD pch_mac l=30n w=100n
MM44_1 net028 SE net030 VDD pch_mac l=30n w=240.00n
MM44_2 net028 SE net030 VDD pch_mac l=30n w=240.00n
MM41 net094 SI VDD VDD pch_mac l=30n w=100n
.ENDS
.SUBCKT SDFQD2 SI D SE CP Q VDD VSS
MM10 net79 qf_x VSS VSS nch_mac l=30.0n w=0.19u
MM9 qf clkb net79 VSS nch_mac l=30.0n w=0.19u
MM27 net124 net68 net0202 VSS nch_mac l=30.0n w=0.175u
MM47 net0202 D VSS VSS nch_mac l=30.0n w=0.175u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.14u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net124 VSS nch_mac l=30.0n w=0.2u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.19u
MM64 mq_x clkbb net111 VSS nch_mac l=30.0n w=0.14u
MM65 net111 mq VSS VSS nch_mac l=30.0n w=0.14u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.19u
MM0 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM2 net124 SE net128 VSS nch_mac l=30.0n w=0.12u
MM3 net128 SI VSS VSS nch_mac l=30.0n w=0.12u
MM14 net68 SE VSS VSS nch_mac l=30.0n w=0.175u
MM6 net8 SI VDD VDD pch_mac l=30.0n w=0.12u
MM7 net12 net68 net8 VDD pch_mac l=30.0n w=0.12u
MM4 qf clkbb net20 VDD pch_mac l=30.0n w=0.18u
MM5 net20 qf_x VDD VDD pch_mac l=30.0n w=0.18u
MM26 net0202 D VDD VDD pch_mac l=30.0n w=0.24u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.18u
MM79 mq_x clkb net35 VDD pch_mac l=30.0n w=0.18u
MM44 net12 SE net0202 VDD pch_mac l=30.0n w=0.24u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.3u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.18u
MM60 net35 mq VDD VDD pch_mac l=30.0n w=0.18u
MM45 mq_x clkbb net12 VDD pch_mac l=30.0n w=0.18u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM1 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM13 net68 SE VDD VDD pch_mac l=30.0n w=0.24u
.ENDS
.SUBCKT SDFQND2 SI D SE CP QN VDD VSS
MM3 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 QN qf VSS VSS nch_mac l=30.0n w=0.14u 
MM10 net76 qf_x VSS VSS nch_mac l=30.0n w=0.12u
MM9 qf clkb net76 VSS nch_mac l=30.0n w=0.12u
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.265u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM64 mq_x clkbb net96 VSS nch_mac l=30.0n w=100n
MM65 net96 mq VSS VSS nch_mac l=30.0n w=100n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.265u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM1 mq_x clkb net132 VSS nch_mac l=30.0n w=0.175u
MM11 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM12 net0232 D VSS VSS nch_mac l=30.0n w=0.175u
MM15 net120 SE VSS VSS nch_mac l=30.0n w=0.175u
MM16 net132 net120 net0232 VSS nch_mac l=30.0n w=0.175u
MM17 net128 SI VSS VSS nch_mac l=30.0n w=0.12u
MM18 net132 SE net128 VSS nch_mac l=30.0n w=0.12u
MM2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM4 qf clkbb net16 VDD pch_mac l=30.0n w=0.285u
MM5 net16 qf_x VDD VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.285u
MM79 mq_x clkb net27 VDD pch_mac l=30.0n w=100n
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.285u
MM60 net27 mq VDD VDD pch_mac l=30.0n w=100n
MM19 net120 SE VDD VDD pch_mac l=30.0n w=0.24u
MM20 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM21 mq_x clkbb net64 VDD pch_mac l=30.0n w=0.2u
MM22 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM23 net64 SE net0232 VDD pch_mac l=30.0n w=0.24u
MM24 net0232 D VDD VDD pch_mac l=30.0n w=0.24u
MM28 net64 net120 net68 VDD pch_mac l=30.0n w=0.12u
MM29 net68 SI VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFQOPTBD2 SI D SE CP Q VDD VSS
MM14 net68 SE VSS VSS nch_mac l=30n w=135.0n
MM3 net088 SI VSS VSS nch_mac l=30n w=100n
MM2 net124 SE net088 VSS nch_mac l=30n w=100n
MM0_1 Q sl_bx VSS VSS nch_mac l=30n w=140.0n
MM0_2 Q sl_bx VSS VSS nch_mac l=30n w=140.0n
MSLTn1 sl_a clkbb ml_b VSS nch_mac l=30n w=220.0n
MM65 net091 ml_b VSS VSS nch_mac l=30n w=100n
MM64 ml_ax clkbb net091 VSS nch_mac l=30n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30n w=130.0n
MM46 ml_ax clkb net124 VSS nch_mac l=30n w=200n
MM76 sl_bx sl_a VSS VSS nch_mac l=30n w=140.0n
MM49_1 ml_b ml_ax VSS VSS nch_mac l=30n w=210.0n
MM49_2 ml_b ml_ax VSS VSS nch_mac l=30n w=210.0n
MM53 clkb CP VSS VSS nch_mac l=30n w=140.0n
MM47_1 net0202 D VSS VSS nch_mac l=30n w=135.0n
MM47_2 net0202 D VSS VSS nch_mac l=30n w=135.0n
MM27_1 net124 net68 net0202 VSS nch_mac l=30n w=210.0n
MM27_2 net124 net68 net0202 VSS nch_mac l=30n w=210.0n
MM9 sl_a clkb net087 VSS nch_mac l=30n w=100n
MM10 net087 sl_bx VSS VSS nch_mac l=30n w=100n
MM17 net0202 D VDD VDD pch_mac l=30n w=170.0n
MM13 net68 SE VDD VDD pch_mac l=30n w=170.0n
MM1_1 Q sl_bx VDD VDD pch_mac l=30n w=170.0n
MM1_2 Q sl_bx VDD VDD pch_mac l=30n w=170.0n
MM8 clkb CP VDD VDD pch_mac l=30n w=170.0n
MM45 ml_ax clkbb net12 VDD pch_mac l=30n w=200n
MM60 net089 ml_b VDD VDD pch_mac l=30n w=100n
MM50_1 ml_b ml_ax VDD VDD pch_mac l=30n w=205.00n
MM50_2 ml_b ml_ax VDD VDD pch_mac l=30n w=205.00n
MM56 clkbb clkb VDD VDD pch_mac l=30n w=300n
MM77 sl_bx sl_a VDD VDD pch_mac l=30n w=170.0n
MM44_1 net12 SE net0202 VDD pch_mac l=30n w=240.00n
MM44_2 net12 SE net0202 VDD pch_mac l=30n w=240.00n
MM79 ml_ax clkb net089 VDD pch_mac l=30n w=100n
MSLTp1 sl_a clkb ml_b VDD pch_mac l=30n w=190.0n
MM26 net0202 D VDD VDD pch_mac l=30n w=170.0n
MM5 net086 sl_bx VDD VDD pch_mac l=30n w=100n
MM4 sl_a clkbb net086 VDD pch_mac l=30n w=100n
MM7 net12 net68 net090 VDD pch_mac l=30n w=100n
MM6 net090 SI VDD VDD pch_mac l=30n w=100n
.ENDS
.SUBCKT SDFSND2 SI D SE CP SDN Q QN VDD VSS
MM32 net86 clkb qf VSS nch_mac l=30.0n w=0.22u
MM7 net86 SDN net93 VSS nch_mac l=30.0n w=0.14u
MM25 mq SDN net98 VSS nch_mac l=30.0n w=0.22u
MM14 net98 mq_x VSS VSS nch_mac l=30.0n w=0.22u
MM9 net93 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM3 QN net86 VSS VSS nch_mac l=30.0n w=0.14u 
MM3_2 QN net86 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM12 net74 D VSS VSS nch_mac l=30.0n w=0.175u
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM64 mq_x clkbb net126 VSS nch_mac l=30.0n w=100n
MM65 net126 mq VSS VSS nch_mac l=30.0n w=100n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.22u
MM11 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM1 mq_x clkb net142 VSS nch_mac l=30.0n w=0.175u
MM18 net142 SE net145 VSS nch_mac l=30.0n w=0.12u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM16 net142 net62 net74 VSS nch_mac l=30.0n w=0.175u
MM17 net145 SI VSS VSS nch_mac l=30.0n w=0.12u
MM15 net62 SE VSS VSS nch_mac l=30.0n w=0.12u
MM2 QN net86 VDD VDD pch_mac l=30.0n w=0.17u 
MM2_2 QN net86 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 net86 qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM30 net86 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM8 net86 SDN VDD VDD pch_mac l=30.0n w=0.12u
MM4 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM10 mq SDN VDD VDD pch_mac l=30.0n w=0.215u
MM13 mq mq_x VDD VDD pch_mac l=30.0n w=0.215u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.31u
MM79 mq_x clkb net45 VDD pch_mac l=30.0n w=100n
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM60 net45 mq VDD VDD pch_mac l=30.0n w=100n
MM20 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM21 mq_x clkbb net78 VDD pch_mac l=30.0n w=0.22u
MM19 net62 SE VDD VDD pch_mac l=30.0n w=0.275u
MM22 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM23 net78 SE net74 VDD pch_mac l=30.0n w=0.275u
MM24 net74 D VDD VDD pch_mac l=30.0n w=0.275u
MM28 net78 net62 net82 VDD pch_mac l=30.0n w=0.12u
MM29 net82 SI VDD VDD pch_mac l=30.0n w=0.12u
.ENDS
.SUBCKT SDFSNQD2 SI D SE CP SDN Q VDD VSS
MM15 net9 SE VSS VSS nch_mac l=30.0n w=0.12u
MM17 net28 SI VSS VSS nch_mac l=30.0n w=0.12u
MM16 net25 net9 net20 VSS nch_mac l=30.0n w=0.175u
MM0 clkbb clkb VSS VSS nch_mac l=30.0n w=0.14u
MM18 net25 SE net28 VSS nch_mac l=30.0n w=0.12u
MM1 mq_x clkb net25 VSS nch_mac l=30.0n w=0.175u
MM11 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.22u
MM65 net48 mq VSS VSS nch_mac l=30.0n w=100n
MM64 mq_x clkbb net48 VSS nch_mac l=30.0n w=100n
MM76 qf_x qf VSS VSS nch_mac l=30.0n w=140.0n
MM12 net20 D VSS VSS nch_mac l=30.0n w=0.175u
MM5 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM9 net76 qf_x VSS VSS nch_mac l=30.0n w=0.14u
MM14 net72 mq_x VSS VSS nch_mac l=30.0n w=0.22u
MM25 mq SDN net72 VSS nch_mac l=30.0n w=0.22u
MM7 net77 SDN net76 VSS nch_mac l=30.0n w=0.14u
MM32 net77 clkb qf VSS nch_mac l=30.0n w=0.22u
MM29 net88 SI VDD VDD pch_mac l=30.0n w=0.12u
MM28 net85 net9 net88 VDD pch_mac l=30.0n w=0.12u
MM24 net20 D VDD VDD pch_mac l=30.0n w=0.275u
MM23 net85 SE net20 VDD pch_mac l=30.0n w=0.275u
MM22 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM19 net9 SE VDD VDD pch_mac l=30.0n w=0.275u
MM21 mq_x clkbb net85 VDD pch_mac l=30.0n w=0.22u
MM20 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM60 net113 mq VDD VDD pch_mac l=30.0n w=100n
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM79 mq_x clkb net113 VDD pch_mac l=30.0n w=100n
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.31u
MM13 mq mq_x VDD VDD pch_mac l=30.0n w=0.215u
MM10 mq SDN VDD VDD pch_mac l=30.0n w=0.215u
MM4 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM8 net77 SDN VDD VDD pch_mac l=30.0n w=0.12u
MM30 net77 clkbb qf VDD pch_mac l=30.0n w=0.12u
MM6 net77 qf_x VDD VDD pch_mac l=30.0n w=170.0n
.ENDS
.SUBCKT SEDFARD2 E SE CP SI D Q QN VDD VSS
MM24 net109 E VSS VSS nch_mac l=30.0n w=0.22u
MM23 net106 D net109 VSS nch_mac l=30.0n w=0.155u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.16u
MM73 QN qf VSS VSS nch_mac l=30.0n w=0.275u 
MM73_2 QN qf VSS VSS nch_mac l=30.0n w=0.275u 
MM48 net157 net174 VSS VSS nch_mac l=30.0n w=140n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.275u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.275u 
MM65 net126 mq_x VSS VSS nch_mac l=30.0n w=0.16u
MM64 mq clkbb net126 VSS nch_mac l=30.0n w=0.16u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=0.29u
MM46 mq clkb net154 VSS nch_mac l=30.0n w=0.16u
MM76 qf qf_x VSS VSS nch_mac l=30.0n w=0.275u
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.16u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=0.29u
MM47 net154 SE net157 VSS nch_mac l=30.0n w=140n
MM20 net106 net86 net161 VSS nch_mac l=30.0n w=0.155u
MM19 net161 qf VSS VSS nch_mac l=30.0n w=0.155u
MM31 qf_x clkb net190 VSS nch_mac l=30.0n w=0.16u
MM16 net170 SE VSS VSS nch_mac l=30.0n w=0.16u
MM14 net174 SI VSS VSS nch_mac l=30.0n w=0.14u
MM28 net178 net170 VSS VSS nch_mac l=30.0n w=0.16u
MM27 net154 net106 net178 VSS nch_mac l=30.0n w=0.14u
MM12 net86 E VSS VSS nch_mac l=30.0n w=0.22u
MM32 net190 qf VSS VSS nch_mac l=30.0n w=0.16u
MM13 net174 SI VDD VDD pch_mac l=30.0n w=0.17u
MM22 net21 net86 VDD VDD pch_mac l=30.0n w=0.25u
MM21 net106 D net21 VDD pch_mac l=30.0n w=0.25u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.31u
MM18 net106 E net30 VDD pch_mac l=30.0n w=0.155u
MM17 net30 qf VDD VDD pch_mac l=30.0n w=0.155u
MM45 mq clkbb net94 VDD pch_mac l=30.0n w=0.205u
MM74 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM74_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM60 net42 mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.31u
MM77 qf qf_x VDD VDD pch_mac l=30.0n w=170n
MM44 net94 net106 net61 VDD pch_mac l=30.0n w=170n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq clkb net42 VDD pch_mac l=30.0n w=0.175u
MM43 net61 SE VDD VDD pch_mac l=30.0n w=0.285u
MM30 net85 qf VDD VDD pch_mac l=30.0n w=0.175u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.175u
MM29 qf_x clkbb net85 VDD pch_mac l=30.0n w=0.175u
MM11 net86 E VDD VDD pch_mac l=30.0n w=0.14u
MM15 net170 SE VDD VDD pch_mac l=30.0n w=0.285u
MM26 net94 net170 net98 VDD pch_mac l=30.0n w=0.17u
MM25 net98 net174 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SEDFCND2 E SE CP SI D CDN Q QN VDD VSS
MM2 net35 net27 net23 VSS nch_mac l=30.0n w=0.14u
MM3 net23 net25 net26 VSS nch_mac l=30.0n w=0.25u
MM0 net27 E VSS VSS nch_mac l=30.0n w=0.275u
MM7 net26 net67 VSS VSS nch_mac l=30.0n w=0.145u
MM52 net35 SE net103 VSS nch_mac l=30.0n w=100n
MM73 net25 qf_x VSS VSS nch_mac l=30.0n w=0.15u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.15u
MM48 net47 E net26 VSS nch_mac l=30.0n w=0.145u
MM67 net25 clkb qf VSS nch_mac l=30.0n w=120.0n
MM69 QN net25 VSS VSS nch_mac l=30.0n w=0.14u 
MM69_2 QN net25 VSS VSS nch_mac l=30.0n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM65 net74 mq net66 VSS nch_mac l=30.0n w=100n
MM57 net67 SE VSS VSS nch_mac l=30.0n w=145.00n
MM64 mq_x clkbb net74 VSS nch_mac l=30.0n w=100n
MM66 net66 CDN VSS VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net35 VSS nch_mac l=30.0n w=0.185u
MM76 qf_x qf net90 VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.26u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM75 net90 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM51 net103 SI VSS VSS nch_mac l=30.0n w=100n
MM47 net35 D net47 VSS nch_mac l=30.0n w=0.14u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
MM1 net27 E VDD VDD pch_mac l=30.0n w=0.12u
MM4 net135 E net131 VDD pch_mac l=30.0n w=0.22u
MM5 net131 net25 net134 VDD pch_mac l=30.0n w=0.22u
MM42 net135 net67 net138 VDD pch_mac l=30.0n w=0.12u
MM6 net134 SE VDD VDD pch_mac l=30.0n w=0.27u
MM45 mq_x clkbb net135 VDD pch_mac l=30.0n w=0.19u
MM70 QN net25 VDD VDD pch_mac l=30.0n w=0.17u 
MM70_2 QN net25 VDD VDD pch_mac l=30.0n w=0.17u 
MM58 net67 SE VDD VDD pch_mac l=30.0n w=135.0n
MM74 net25 qf_x VDD VDD pch_mac l=30.0n w=0.275u
MM60 net159 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM41 net138 SI VDD VDD pch_mac l=30.0n w=0.12u
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.22u
MM61 net159 mq VDD VDD pch_mac l=30.0n w=120.0n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=275.00n
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM44 net135 D net190 VDD pch_mac l=30.0n w=0.22u
MM68 net25 clkbb qf VDD pch_mac l=30.0n w=275.00n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq_x clkb net159 VDD pch_mac l=30.0n w=0.12u
MM43 net190 net27 net134 VDD pch_mac l=30.0n w=0.22u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
.ENDS
.SUBCKT SEDFCNQD2 E SE CP SI D CDN Q VDD VSS
MM47 net166 D net154 VSS nch_mac l=30.0n w=0.14u
MM51 net169 SI VSS VSS nch_mac l=30.0n w=100n
MM75 net106 CDN VSS VSS nch_mac l=30.0n w=140.0n
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq mq_x VSS VSS nch_mac l=30.0n w=0.26u
MM76 qf_x qf net106 VSS nch_mac l=30.0n w=140.0n
MM46 mq_x clkb net166 VSS nch_mac l=30.0n w=0.185u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM66 net130 CDN VSS VSS nch_mac l=30.0n w=100n
MM64 mq_x clkbb net137 VSS nch_mac l=30.0n w=100n
MM57 net138 SE VSS VSS nch_mac l=30.0n w=145.00n
MM65 net137 mq net130 VSS nch_mac l=30.0n w=100n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM67 net180 clkb qf VSS nch_mac l=30.0n w=120.0n
MM48 net154 E net181 VSS nch_mac l=30.0n w=0.145u
MSLTn1 qf clkbb mq VSS nch_mac l=30.0n w=0.15u
MM73 net180 qf_x VSS VSS nch_mac l=30.0n w=0.15u
MM52 net166 SE net169 VSS nch_mac l=30.0n w=100n
MM7 net181 net138 VSS VSS nch_mac l=30.0n w=0.145u
MM0 net90 E VSS VSS nch_mac l=30.0n w=0.275u
MM3 net185 net180 net181 VSS nch_mac l=30.0n w=0.25u
MM2 net166 net90 net185 VSS nch_mac l=30.0n w=0.14u
MSLTp1 qf clkb mq VDD pch_mac l=30.0n w=0.275u
MM43 net14 net90 net85 VDD pch_mac l=30.0n w=0.22u
MM79 mq_x clkb net21 VDD pch_mac l=30.0n w=0.12u
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM68 net180 clkbb qf VDD pch_mac l=30.0n w=275.00n
MM44 net78 D net14 VDD pch_mac l=30.0n w=0.22u
MM77 qf_x qf VDD VDD pch_mac l=30.0n w=170.0n
MM78 qf_x CDN VDD VDD pch_mac l=30.0n w=275.00n
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.17u
MM61 net21 mq VDD VDD pch_mac l=30.0n w=120.0n
MM50 mq mq_x VDD VDD pch_mac l=30.0n w=0.22u
MM41 net81 SI VDD VDD pch_mac l=30.0n w=0.12u
MM60 net21 CDN VDD VDD pch_mac l=30.0n w=0.12u
MM74 net180 qf_x VDD VDD pch_mac l=30.0n w=0.275u
MM58 net138 SE VDD VDD pch_mac l=30.0n w=135.0n
MM45 mq_x clkbb net78 VDD pch_mac l=30.0n w=0.19u
MM6 net85 SE VDD VDD pch_mac l=30.0n w=0.27u
MM42 net78 net138 net81 VDD pch_mac l=30.0n w=0.12u
MM5 net82 net180 net85 VDD pch_mac l=30.0n w=0.22u
MM4 net78 E net82 VDD pch_mac l=30.0n w=0.22u
MM1 net90 E VDD VDD pch_mac l=30.0n w=0.12u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SEDFD2 E SE CP SI D Q QN VDD VSS
MM24 net109 E VSS VSS nch_mac l=30.0n w=0.22u
MM23 net106 D net109 VSS nch_mac l=30.0n w=0.155u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.26u
MM73 QN qf VSS VSS nch_mac l=30.0n w=0.275u 
MM73_2 QN qf VSS VSS nch_mac l=30.0n w=0.275u 
MM48 net157 net174 VSS VSS nch_mac l=30.0n w=140.0n
MM71 Q qf_x VSS VSS nch_mac l=30.0n w=0.275u 
MM71_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.275u 
MM65 net126 mq_x VSS VSS nch_mac l=30.0n w=100n
MM64 mq clkbb net126 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq clkb net154 VSS nch_mac l=30.0n w=190.0n
MM76 qf qf_x VSS VSS nch_mac l=30.0n w=0.275u
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM47 net154 SE net157 VSS nch_mac l=30.0n w=140.0n
MM20 net106 net86 net161 VSS nch_mac l=30.0n w=0.155u
MM19 net161 qf VSS VSS nch_mac l=30.0n w=0.155u
MM31 qf_x clkb net190 VSS nch_mac l=30.0n w=0.12u
MM16 net170 SE VSS VSS nch_mac l=30.0n w=0.16u
MM14 net174 SI VSS VSS nch_mac l=30.0n w=0.14u
MM28 net178 net170 VSS VSS nch_mac l=30.0n w=0.16u
MM27 net154 net106 net178 VSS nch_mac l=30.0n w=0.14u
MM12 net86 E VSS VSS nch_mac l=30.0n w=0.22u
MM32 net190 qf VSS VSS nch_mac l=30.0n w=0.12u
MM13 net174 SI VDD VDD pch_mac l=30.0n w=0.17u
MM22 net21 net86 VDD VDD pch_mac l=30.0n w=0.25u
MM21 net106 D net21 VDD pch_mac l=30.0n w=0.25u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.33u
MM18 net106 E net30 VDD pch_mac l=30.0n w=0.155u
MM17 net30 qf VDD VDD pch_mac l=30.0n w=0.155u
MM45 mq clkbb net94 VDD pch_mac l=30.0n w=200n
MM74 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM74_2 QN qf VDD VDD pch_mac l=30.0n w=0.17u 
MM60 net42 mq_x VDD VDD pch_mac l=30.0n w=100n
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.295u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.33u
MM77 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM44 net94 net106 net61 VDD pch_mac l=30.0n w=170.0n
MM72 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM79 mq clkb net42 VDD pch_mac l=30.0n w=100n
MM43 net61 SE VDD VDD pch_mac l=30.0n w=0.285u
MM30 net85 qf VDD VDD pch_mac l=30.0n w=0.12u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.295u
MM29 qf_x clkbb net85 VDD pch_mac l=30.0n w=0.295u
MM11 net86 E VDD VDD pch_mac l=30.0n w=0.12u
MM15 net170 SE VDD VDD pch_mac l=30.0n w=0.285u
MM26 net94 net170 net98 VDD pch_mac l=30.0n w=0.17u
MM25 net98 net174 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT SEDFQARD2 E SE CP SI D Q VDD VSS
MM0 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM2 net101 SE VSS VSS nch_mac l=30.0n w=0.16u
MM24 net24 E VSS VSS nch_mac l=30.0n w=0.22u
MM23 net21 D net24 VSS nch_mac l=30.0n w=0.155u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.16u
MM48 net29 net165 VSS VSS nch_mac l=30.0n w=140n
MM65 net40 mq_x VSS VSS nch_mac l=30.0n w=0.16u
MM64 mq clkbb net40 VSS nch_mac l=30.0n w=0.16u
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140n
MM46 mq clkb net61 VSS nch_mac l=30.0n w=0.16u
MM76 qf qf_x VSS VSS nch_mac l=30.0n w=140n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.16u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140n
MM47 net61 SE net29 VSS nch_mac l=30.0n w=140n
MM20 net21 net120 net69 VSS nch_mac l=30.0n w=0.155u
MM19 net69 qf VSS VSS nch_mac l=30.0n w=0.155u
MM16 net165 SI VSS VSS nch_mac l=30.0n w=0.14u
MM14 net120 E VSS VSS nch_mac l=30.0n w=0.22u
MM28 net81 net101 VSS VSS nch_mac l=30.0n w=0.16u
MM27 net61 net21 net81 VSS nch_mac l=30.0n w=0.14u
MM9 qf_x clkb net93 VSS nch_mac l=30.0n w=0.16u
MM10 net93 qf VSS VSS nch_mac l=30.0n w=0.16u
MM1 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net101 SE VDD VDD pch_mac l=30.0n w=0.285u
MM13 net120 E VDD VDD pch_mac l=30.0n w=0.14u
MM22 net116 net120 VDD VDD pch_mac l=30.0n w=0.25u
MM21 net21 D net116 VDD pch_mac l=30.0n w=0.25u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.33u
MM18 net21 E net125 VDD pch_mac l=30.0n w=0.155u
MM17 net125 qf VDD VDD pch_mac l=30.0n w=0.155u
MM45 mq clkbb net169 VDD pch_mac l=30.0n w=0.205u
MM60 net156 mq_x VDD VDD pch_mac l=30.0n w=0.175u
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.175u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.33u
MM77 qf qf_x VDD VDD pch_mac l=30.0n w=170n
MM44 net169 net21 net157 VDD pch_mac l=30.0n w=170n
MM79 mq clkb net156 VDD pch_mac l=30.0n w=0.175u
MM43 net157 SE VDD VDD pch_mac l=30.0n w=0.285u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.175u
MM15 net165 SI VDD VDD pch_mac l=30.0n w=0.17u
MM26 net169 net101 net172 VDD pch_mac l=30.0n w=0.17u
MM25 net172 net165 VDD VDD pch_mac l=30.0n w=0.17u
MM5 net177 qf VDD VDD pch_mac l=30.0n w=0.175u
MM4 qf_x clkbb net177 VDD pch_mac l=30.0n w=0.175u
.ENDS
.SUBCKT SEDFQD2 E SE CP SI D Q VDD VSS
MM0 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Q qf_x VSS VSS nch_mac l=30.0n w=0.14u 
MM2 net101 SE VSS VSS nch_mac l=30.0n w=0.16u
MM24 net24 E VSS VSS nch_mac l=30.0n w=0.22u
MM23 net21 D net24 VSS nch_mac l=30.0n w=0.155u
MSLTn1 qf_x clkbb mq_x VSS nch_mac l=30.0n w=0.26u
MM48 net29 net165 VSS VSS nch_mac l=30.0n w=140.0n
MM65 net40 mq_x VSS VSS nch_mac l=30.0n w=100n
MM64 mq clkbb net40 VSS nch_mac l=30.0n w=100n
MM55 clkbb clkb VSS VSS nch_mac l=30.0n w=140.0n
MM46 mq clkb net61 VSS nch_mac l=30.0n w=190.0n
MM76 qf qf_x VSS VSS nch_mac l=30.0n w=140.0n
MM49 mq_x mq VSS VSS nch_mac l=30.0n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30.0n w=140.0n
MM47 net61 SE net29 VSS nch_mac l=30.0n w=140.0n
MM20 net21 net120 net69 VSS nch_mac l=30.0n w=0.155u
MM19 net69 qf VSS VSS nch_mac l=30.0n w=0.155u
MM16 net165 SI VSS VSS nch_mac l=30.0n w=0.14u
MM14 net120 E VSS VSS nch_mac l=30.0n w=0.22u
MM28 net81 net101 VSS VSS nch_mac l=30.0n w=0.16u
MM27 net61 net21 net81 VSS nch_mac l=30.0n w=0.14u
MM9 qf_x clkb net93 VSS nch_mac l=30.0n w=0.12u
MM10 net93 qf VSS VSS nch_mac l=30.0n w=0.12u
MM1 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Q qf_x VDD VDD pch_mac l=30.0n w=0.17u 
MM3 net101 SE VDD VDD pch_mac l=30.0n w=0.285u
MM13 net120 E VDD VDD pch_mac l=30.0n w=0.12u
MM22 net116 net120 VDD VDD pch_mac l=30.0n w=0.25u
MM21 net21 D net116 VDD pch_mac l=30.0n w=0.25u
MM8 clkb CP VDD VDD pch_mac l=30.0n w=0.33u
MM18 net21 E net125 VDD pch_mac l=30.0n w=0.155u
MM17 net125 qf VDD VDD pch_mac l=30.0n w=0.155u
MM45 mq clkbb net169 VDD pch_mac l=30.0n w=200n
MM60 net156 mq_x VDD VDD pch_mac l=30.0n w=100n
MM50 mq_x mq VDD VDD pch_mac l=30.0n w=0.295u
MM56 clkbb clkb VDD VDD pch_mac l=30.0n w=0.33u
MM77 qf qf_x VDD VDD pch_mac l=30.0n w=170.0n
MM44 net169 net21 net157 VDD pch_mac l=30.0n w=170.0n
MM79 mq clkb net156 VDD pch_mac l=30.0n w=100n
MM43 net157 SE VDD VDD pch_mac l=30.0n w=0.285u
MSLTp1 qf_x clkb mq_x VDD pch_mac l=30.0n w=0.295u
MM15 net165 SI VDD VDD pch_mac l=30.0n w=0.17u
MM26 net169 net101 net172 VDD pch_mac l=30.0n w=0.17u
MM25 net172 net165 VDD VDD pch_mac l=30.0n w=0.17u
MM5 net177 qf VDD VDD pch_mac l=30.0n w=0.12u
MM4 qf_x clkbb net177 VDD pch_mac l=30.0n w=0.295u
.ENDS
.SUBCKT XNR2D2 A1 A2 ZN VDD VSS
MM6 ZN net093 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 ZN net093 VSS VSS nch_mac l=30.0n w=0.14u 
MM8 net17 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM17 net26 A1 net093 VSS nch_mac l=30.0n w=0.205u
MM3 net46 net17 net093 VSS nch_mac l=30.0n w=0.205u
MM5 net46 net26 VSS VSS nch_mac l=30.0n w=0.14u
MM0 net26 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM7 ZN net093 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 ZN net093 VDD VDD pch_mac l=30.0n w=0.17u 
MM9 net17 A1 VDD VDD pch_mac l=30.0n w=0.33u
MM16 net26 net17 net093 VDD pch_mac l=30.0n w=0.17u
MM4 net46 A1 net093 VDD pch_mac l=30.0n w=0.17u
MM1 net46 net26 VDD VDD pch_mac l=30.0n w=0.33u
MM2 net26 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT XNR2OPTND2 A1 A2 ZN VDD VSS
MM0_1 net3 A2 VDD VDD pch_mac l=30n w=170.0n
MM0_2 net3 A2 VDD VDD pch_mac l=30n w=170.0n
MM3_1 net7 net3 VDD VDD pch_mac l=30n w=170.0n
MM3_2 net7 net3 VDD VDD pch_mac l=30n w=170.0n
MM4_1 ZN net15 net7 VDD pch_mac l=30n w=170.0n
MM4_2 ZN net15 net7 VDD pch_mac l=30n w=170.0n
MM7_1 ZN A1 net3 VDD pch_mac l=30n w=170.0n
MM7_2 ZN A1 net3 VDD pch_mac l=30n w=170.0n
MM9 net15 A1 VDD VDD pch_mac l=30n w=170.0n
MM1_1 net3 A2 VSS VSS nch_mac l=30n w=140.0n
MM1_2 net3 A2 VSS VSS nch_mac l=30n w=140.0n
MM2_1 net7 net3 VSS VSS nch_mac l=30n w=140.0n
MM2_2 net7 net3 VSS VSS nch_mac l=30n w=140.0n
MM5_1 ZN A1 net7 VSS nch_mac l=30n w=140.0n
MM5_2 ZN A1 net7 VSS nch_mac l=30n w=140.0n
MM6_1 ZN net15 net3 VSS nch_mac l=30n w=140.0n
MM6_2 ZN net15 net3 VSS nch_mac l=30n w=140.0n
MM8 net15 A1 VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT XNR3D2 A1 A2 A3 ZN VDD VSS
MM5 net082 net179 VSS VSS nch_mac l=30.0n w=0.205u
MM7 net082 net191 net230 VSS nch_mac l=30.0n w=0.205u
MM19 net195 net187 VSS VSS nch_mac l=30.0n w=140.0n
MM18 net195 net211 net206 VSS nch_mac l=30.0n w=140.0n
MM8 net191 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM0 net187 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM17 net179 A2 net230 VSS nch_mac l=30.0n w=0.205u
MM3 net179 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM11 net187 net230 net206 VSS nch_mac l=30.0n w=140.0n
MM13 net211 net230 VSS VSS nch_mac l=30.0n w=0.14u
MM21 ZN net206 VSS VSS nch_mac l=30.0n w=0.14u 
MM21_2 ZN net206 VSS VSS nch_mac l=30.0n w=0.14u 
MM14 net195 net230 net206 VDD pch_mac l=30.0n w=0.265u
MM15 net195 net187 VDD VDD pch_mac l=30.0n w=0.315u
MM6 net082 A2 net230 VDD pch_mac l=30.0n w=0.275u
MM20 ZN net206 VDD VDD pch_mac l=30.0n w=0.17u 
MM20_2 ZN net206 VDD VDD pch_mac l=30.0n w=0.17u 
MM4 net082 net179 VDD VDD pch_mac l=30.0n w=0.21u
MM9 net191 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM2 net187 A3 VDD VDD pch_mac l=30.0n w=0.17u
MM16 net179 net191 net230 VDD pch_mac l=30.0n w=0.275u
MM1 net179 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM10 net187 net211 net206 VDD pch_mac l=30.0n w=0.265u
MM12 net211 net230 VDD VDD pch_mac l=30.0n w=0.315u
.ENDS
.SUBCKT XNR4D2 A1 A2 A3 A4 ZN VDD VSS
MM4 net16 net124 VSS VSS nch_mac l=30.0n w=0.14u
MM5 net16 A1 net71 VSS nch_mac l=30.0n w=0.14u
MM43 ZN net91 VSS VSS nch_mac l=30.0n w=0.14u 
MM43_2 ZN net91 VSS VSS nch_mac l=30.0n w=0.14u 
MM41 net36 net0187 net91 VSS nch_mac l=30.0n w=0.14u
MM40 net71 net107 net91 VSS nch_mac l=30.0n w=0.14u
MM37 net107 net0187 VSS VSS nch_mac l=30.0n w=140.0n
MM35 net36 net71 VSS VSS nch_mac l=30.0n w=0.14u
MM31 net0180 A4 VSS VSS nch_mac l=30.0n w=0.14u
MM27 net116 net0180 net0187 VSS nch_mac l=30.0n w=0.14u
MM29 net48 net116 VSS VSS nch_mac l=30.0n w=0.14u
MM28 net48 A4 net0187 VSS nch_mac l=30.0n w=0.14u
MM30 net116 A3 VSS VSS nch_mac l=30.0n w=140.0n
MM17 net124 net60 net71 VSS nch_mac l=30.0n w=0.14u
MM8 net60 A1 VSS VSS nch_mac l=30.0n w=140.0n
MM3 net124 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM2 net16 net60 net71 VDD pch_mac l=30.0n w=0.17u
MM0 net16 net124 VDD VDD pch_mac l=30.0n w=0.27u
MM42 ZN net91 VDD VDD pch_mac l=30.0n w=0.17u 
MM42_2 ZN net91 VDD VDD pch_mac l=30.0n w=0.17u 
MM39 net36 net107 net91 VDD pch_mac l=30.0n w=0.17u
MM38 net71 net0187 net91 VDD pch_mac l=30.0n w=0.17u
MM36 net107 net0187 VDD VDD pch_mac l=30.0n w=170.0n
MM34 net36 net71 VDD VDD pch_mac l=30.0n w=0.17u
MM26 net0180 A4 VDD VDD pch_mac l=30.0n w=0.17u
MM22 net116 A4 net0187 VDD pch_mac l=30.0n w=0.17u
MM24 net48 net116 VDD VDD pch_mac l=30.0n w=0.17u
MM23 net48 net0180 net0187 VDD pch_mac l=30.0n w=0.17u
MM25 net116 A3 VDD VDD pch_mac l=30.0n w=170.0n
MM16 net124 A1 net71 VDD pch_mac l=30.0n w=0.17u
MM9 net60 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM1 net124 A2 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT XOR2D2 A1 A2 Z VDD VSS
MM3 net10 A1 net14 VSS nch_mac l=30.0n w=0.205u
MM17 net10 net36 net13 VSS nch_mac l=30.0n w=0.205u
MM5 net14 net13 VSS VSS nch_mac l=30.0n w=0.245u
MM6 Z net10 VSS VSS nch_mac l=30.0n w=0.14u 
MM6_2 Z net10 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net13 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net36 A1 VSS VSS nch_mac l=30.0n w=0.245u
MM16 net10 A1 net13 VDD pch_mac l=30.0n w=0.17u
MM1 net14 net13 VDD VDD pch_mac l=30.0n w=0.245u
MM2 net13 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM9 net36 A1 VDD VDD pch_mac l=30.0n w=0.245u
MM7 Z net10 VDD VDD pch_mac l=30.0n w=0.17u 
MM7_2 Z net10 VDD VDD pch_mac l=30.0n w=0.17u 
MM4 net10 net36 net14 VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT XOR2OPTND2 A1 A2 Z VDD VSS
MM0_1 net3 A2 VDD VDD pch_mac l=30n w=170.0n
MM0_2 net3 A2 VDD VDD pch_mac l=30n w=170.0n
MM3_1 net7 net3 VDD VDD pch_mac l=30n w=170.0n
MM3_2 net7 net3 VDD VDD pch_mac l=30n w=170.0n
MM4_1 Z A1 net7 VDD pch_mac l=30n w=170.0n
MM4_2 Z A1 net7 VDD pch_mac l=30n w=170.0n
MM7_1 Z net15 net3 VDD pch_mac l=30n w=170.0n
MM7_2 Z net15 net3 VDD pch_mac l=30n w=170.0n
MM9 net15 A1 VDD VDD pch_mac l=30n w=170.0n
MM1_1 net3 A2 VSS VSS nch_mac l=30n w=140.0n
MM1_2 net3 A2 VSS VSS nch_mac l=30n w=140.0n
MM2_1 net7 net3 VSS VSS nch_mac l=30n w=140.0n
MM2_2 net7 net3 VSS VSS nch_mac l=30n w=140.0n
MM5_1 Z net15 net7 VSS nch_mac l=30n w=140.0n
MM5_2 Z net15 net7 VSS nch_mac l=30n w=140.0n
MM6_1 Z A1 net3 VSS nch_mac l=30n w=140.0n
MM6_2 Z A1 net3 VSS nch_mac l=30n w=140.0n
MM8 net15 A1 VSS VSS nch_mac l=30n w=140.0n
.ENDS
.SUBCKT XOR3D2 A1 A2 A3 Z VDD VSS
MM21 Z net18 VSS VSS nch_mac l=30.0n w=0.14u 
MM21_2 Z net18 VSS VSS nch_mac l=30.0n w=0.14u 
MM13 net11 net63 VSS VSS nch_mac l=30.0n w=0.14u
MM11 net27 net63 net18 VSS nch_mac l=30.0n w=140.0n
MM3 net19 A1 VSS VSS nch_mac l=30.0n w=0.14u
MM17 net63 net31 net19 VSS nch_mac l=30.0n w=275.00n
MM0 net27 A3 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net31 A2 VSS VSS nch_mac l=30.0n w=140.0n
MM18 net87 net11 net18 VSS nch_mac l=30.0n w=140.0n
MM19 net87 net27 VSS VSS nch_mac l=30.0n w=140.0n
MM7 net0167 A2 net63 VSS nch_mac l=30.0n w=275.00n
MM5 net0167 net19 VSS VSS nch_mac l=30.0n w=275.00n
MM12 net11 net63 VDD VDD pch_mac l=30.0n w=0.315u
MM10 net27 net11 net18 VDD pch_mac l=30.0n w=0.265u
MM1 net19 A1 VDD VDD pch_mac l=30.0n w=0.17u
MM16 net63 A2 net19 VDD pch_mac l=30.0n w=0.275u
MM2 net27 A3 VDD VDD pch_mac l=30.0n w=0.17u
MM9 net31 A2 VDD VDD pch_mac l=30.0n w=170.0n
MM4 net0167 net19 VDD VDD pch_mac l=30.0n w=0.33u
MM20 Z net18 VDD VDD pch_mac l=30.0n w=0.17u 
MM20_2 Z net18 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 net0167 net31 net63 VDD pch_mac l=30.0n w=0.275u
MM15 net87 net27 VDD VDD pch_mac l=30.0n w=0.315u
MM14 net87 net63 net18 VDD pch_mac l=30.0n w=0.265u
.ENDS
.SUBCKT XOR4D2 A1 A2 A3 A4 Z VDD VSS
MM3 net8 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net12 A1 VSS VSS nch_mac l=30.0n w=140.0n
MM17 net8 net12 net19 VSS nch_mac l=30.0n w=275.00n
MM30 net80 A3 VSS VSS nch_mac l=30.0n w=140.0n
MM28 net88 A4 net0120 VSS nch_mac l=30.0n w=150.0n
MM29 net88 net80 VSS VSS nch_mac l=30.0n w=150.0n
MM27 net80 net0181 net0120 VSS nch_mac l=30.0n w=150.0n
MM31 net0181 A4 VSS VSS nch_mac l=30.0n w=150.0n
MM35 net100 net19 VSS VSS nch_mac l=30.0n w=0.2u
MM37 net35 net0120 VSS VSS nch_mac l=30.0n w=0.2u
MM40 net19 net0120 net51 VSS nch_mac l=30.0n w=0.16u
MM41 net100 net35 net51 VSS nch_mac l=30.0n w=0.16u
MM43 Z net51 VSS VSS nch_mac l=30.0n w=0.14u 
MM43_2 Z net51 VSS VSS nch_mac l=30.0n w=0.14u 
MM5 net64 A1 net19 VSS nch_mac l=30.0n w=275.00n
MM4 net64 net8 VSS VSS nch_mac l=30.0n w=275.00n
MM1 net8 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM9 net12 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM16 net8 A1 net19 VDD pch_mac l=30.0n w=0.26u
MM25 net80 A3 VDD VDD pch_mac l=30.0n w=170.0n
MM23 net88 net0181 net0120 VDD pch_mac l=30.0n w=165.00n
MM24 net88 net80 VDD VDD pch_mac l=30.0n w=170.0n
MM22 net80 A4 net0120 VDD pch_mac l=30.0n w=165.00n
MM26 net0181 A4 VDD VDD pch_mac l=30.0n w=0.17u
MM34 net100 net19 VDD VDD pch_mac l=30.0n w=0.17u
MM36 net35 net0120 VDD VDD pch_mac l=30.0n w=0.17u
MM38 net19 net35 net51 VDD pch_mac l=30.0n w=0.165u
MM39 net100 net0120 net51 VDD pch_mac l=30.0n w=0.165u
MM42 Z net51 VDD VDD pch_mac l=30.0n w=0.17u 
MM42_2 Z net51 VDD VDD pch_mac l=30.0n w=0.17u 
MM0 net64 net8 VDD VDD pch_mac l=30.0n w=170.0n
MM2 net64 net12 net19 VDD pch_mac l=30.0n w=0.26u
.ENDS
.SUBCKT SDFNSYNCND2 SI D SE CPN CDN Q QN VDD VSS
MM6 qf clkb net0154 VSS nch_mac l=30n w=0.14u
MM7 net0154 net0232 VSS VSS nch_mac l=30n w=0.14u
MM12 net0171 SE net0172 VSS nch_mac l=30n w=0.12u
MM27 net0171 D net0187 VSS nch_mac l=30n w=0.22u
MM14 net0183 SE VSS VSS nch_mac l=30n w=0.22u
MM0 net0232 net0301 VSS VSS nch_mac l=30n w=0.14u
MM2 net0200 net0232 VSS VSS nch_mac l=30n w=0.14u
MM11 net0172 SI VSS VSS nch_mac l=30n w=0.12u
MM26 net0156 CDN net0148 VSS nch_mac l=30n w=0.14u
MM46 mq_x clkbb net0171 VSS nch_mac l=30n w=0.14u
MM47 net0187 net0183 VSS VSS nch_mac l=30n w=0.22u
MM28 mq_x clkb net0156 VSS nch_mac l=30n w=0.14u
MM73 net102 qf_x VSS VSS nch_mac l=30n w=0.14u
MM23 net102 clkbb qf VSS nch_mac l=30n w=0.14u
MM69 QN net102 VSS VSS nch_mac l=30n w=0.14u 
MM69_2 QN net102 VSS VSS nch_mac l=30n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM29 net0148 net0200 VSS VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM76 qf_x qf net150 VSS nch_mac l=30n w=0.14u
MM49 net0301 mq_x VSS VSS nch_mac l=30n w=0.14u
MM53 clkb CPN VSS VSS nch_mac l=30n w=0.14u
MM75 net150 CDN VSS VSS nch_mac l=30n w=0.14u
MM3 net0200 net0232 VDD VDD pch_mac l=30n w=0.17u
MM9 qf clkbb net0236 VDD pch_mac l=30n w=0.17u
MM10 net0236 net0232 VDD VDD pch_mac l=30n w=0.17u
MM1 net0232 net0301 VDD VDD pch_mac l=30n w=0.17u
MM70 QN net102 VDD VDD pch_mac l=30n w=0.335u 
MM70_2 QN net102 VDD VDD pch_mac l=30n w=0.335u 
MM74 net102 qf_x VDD VDD pch_mac l=30n w=0.335u
MM5 net0234 CDN VDD VDD pch_mac l=30n w=0.17u
MM50 net0301 mq_x VDD VDD pch_mac l=30n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM13 net102 clkb qf VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM54 clkb CPN VDD VDD pch_mac l=30n w=0.17u
MM16 net0183 SE VDD VDD pch_mac l=30n w=0.21u
MM45 mq_x clkb net0262 VDD pch_mac l=30n w=0.17u
MM44 net0262 D net0266 VDD pch_mac l=30n w=0.21u
MM15 mq_x clkbb net0234 VDD pch_mac l=30n w=0.17u
MM8 net0234 net0200 VDD VDD pch_mac l=30n w=0.17u
MM17 net0266 SE VDD VDD pch_mac l=30n w=0.21u
MM18 net0262 net0183 net0258 VDD pch_mac l=30n w=100n
MM19 net0258 SI VDD VDD pch_mac l=30n w=100n
.ENDS
.SUBCKT SDFNSYNCSND2 SI D SE CPN CDN SDN Q QN VDD VSS
MM21 net18 net23 VDD VDD pch_mac l=30n w=0.17u
MM16 net167 net23 VDD VDD pch_mac l=30n w=0.17u
MM15 net23 mq VDD VDD pch_mac l=30n w=0.17u
MM20 qf clkbb net18 VDD pch_mac l=30n w=0.17u
MM1 mq net59 VDD VDD pch_mac l=30n w=0.17u
MM54 clkb CPN VDD VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM43 net90 SE VDD VDD pch_mac l=30n w=0.21u
MM11 net91 CDN VDD VDD pch_mac l=30n w=0.17u
MM14 net132 clkb qf VDD pch_mac l=30n w=0.17u
MM44 net55 D net90 VDD pch_mac l=30n w=0.21u
MM77 qf_x CDN VDD VDD pch_mac l=30n w=0.33u
MM78 qf_x qf VDD VDD pch_mac l=30n w=0.33u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM12 net59 clkbb net91 VDD pch_mac l=30n w=0.17u
MM0 mq SDN VDD VDD pch_mac l=30n w=0.17u
MM41 net58 SI VDD VDD pch_mac l=30n w=0.12u
MM13 net91 net167 VDD VDD pch_mac l=30n w=0.17u
MM58 net172 SE VDD VDD pch_mac l=30n w=0.21u
MM70 QN net132 VDD VDD pch_mac l=30n w=0.17u 
MM70_2 QN net132 VDD VDD pch_mac l=30n w=0.17u 
MM45 net59 clkb net55 VDD pch_mac l=30n w=0.17u
MM42 net55 net172 net58 VDD pch_mac l=30n w=0.12u
MM4 net132 qf_x VDD VDD pch_mac l=30n w=0.33u
MM5 net132 SDN VDD VDD pch_mac l=30n w=0.33u
MM18 qf clkb net108 VSS nch_mac l=30n w=0.14u
MM49 net23 mq VSS VSS nch_mac l=30n w=0.14u
MM17 net167 net23 VSS VSS nch_mac l=30n w=0.14u
MM19 net108 net23 VSS VSS nch_mac l=30n w=0.14u
MM75 net145 qf VSS VSS nch_mac l=30n w=0.275u
MM47 net160 D net164 VSS nch_mac l=30n w=0.22u
MM51 net161 SI VSS VSS nch_mac l=30n w=0.12u
MM46 net59 clkbb net160 VSS nch_mac l=30n w=0.14u
MM53 clkb CPN VSS VSS nch_mac l=30n w=0.14u
MM76 qf_x CDN net145 VSS nch_mac l=30n w=0.275u
MM9 net59 clkb net177 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.135u
MM8 net177 CDN net181 VSS nch_mac l=30n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM57 net172 SE VSS VSS nch_mac l=30n w=0.22u
MM10 net181 net167 VSS VSS nch_mac l=30n w=0.14u
MM48 net164 net172 VSS VSS nch_mac l=30n w=0.22u
MM69 QN net132 VSS VSS nch_mac l=30n w=0.14u 
MM69_2 QN net132 VSS VSS nch_mac l=30n w=0.14u 
MM50 net132 clkbb qf VSS nch_mac l=30n w=0.14u
MM2 mq SDN net157 VSS nch_mac l=30n w=0.14u
MM52 net160 SE net161 VSS nch_mac l=30n w=0.12u
MM6 net132 SDN net125 VSS nch_mac l=30n w=0.275u
MM3 net157 net59 VSS VSS nch_mac l=30n w=0.14u
MM7 net125 qf_x VSS VSS nch_mac l=30n w=0.275u
.ENDS
.SUBCKT SDFNSYND2 SI D SE CPN Q QN VDD VSS
MM0 net243 net275 VSS VSS nch_mac l=30n w=0.14u
MM5 net183 net243 VSS VSS nch_mac l=30n w=0.14u
MM47 net211 D net203 VSS nch_mac l=30n w=0.22u
MM51 net214 SI VSS VSS nch_mac l=30n w=0.12u
MM53 clkb CPN VSS VSS nch_mac l=30n w=0.14u
MM49 net275 mq_x VSS VSS nch_mac l=30n w=0.14u
MM46 mq_x clkbb net211 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM26 net193 net183 VSS VSS nch_mac l=30n w=0.14u
MM57 net283 SE VSS VSS nch_mac l=30n w=0.22u
MM28 mq_x clkb net193 VSS nch_mac l=30n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM30 net200 clkbb qf VSS nch_mac l=30n w=0.14u
MM48 net203 net283 VSS VSS nch_mac l=30n w=0.22u
MM7 net208 net243 VSS VSS nch_mac l=30n w=0.14u
MM52 net211 SE net214 VSS nch_mac l=30n w=0.12u
MM2 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM69 QN net200 VSS VSS nch_mac l=30n w=0.14u 
MM69_2 QN net200 VSS VSS nch_mac l=30n w=0.14u 
MM73 net200 qf_x VSS VSS nch_mac l=30n w=0.14u
MM9 qf clkb net208 VSS nch_mac l=30n w=0.14u
MM4 net183 net243 VDD VDD pch_mac l=30n w=0.17u
MM12 net235 net243 VDD VDD pch_mac l=30n w=0.17u
MM13 qf clkbb net235 VDD pch_mac l=30n w=0.17u
MM3 net243 net275 VDD VDD pch_mac l=30n w=0.17u
MM54 clkb CPN VDD VDD pch_mac l=30n w=0.17u
MM43 net251 SE VDD VDD pch_mac l=30n w=0.21u
MM6 net298 net183 VDD VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM8 net200 clkb qf VDD pch_mac l=30n w=0.17u
MM44 net291 D net251 VDD pch_mac l=30n w=0.21u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM50 net275 mq_x VDD VDD pch_mac l=30n w=0.17u
MM41 net279 SI VDD VDD pch_mac l=30n w=100n
MM58 net283 SE VDD VDD pch_mac l=30n w=0.21u
MM45 mq_x clkb net291 VDD pch_mac l=30n w=0.17u
MM42 net291 net283 net279 VDD pch_mac l=30n w=100n
MM16 mq_x clkbb net298 VDD pch_mac l=30n w=0.17u
MM1 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM74 net200 qf_x VDD VDD pch_mac l=30n w=0.17u
MM70 QN net200 VDD VDD pch_mac l=30n w=0.17u 
MM70_2 QN net200 VDD VDD pch_mac l=30n w=0.17u 
.ENDS
.SUBCKT SDFNSYNSND2 SI D SE CPN SDN Q QN VDD VSS
MM35 net10 net111 VDD VDD pch_mac l=30n w=0.17u
MM34 qf clkbb net10 VDD pch_mac l=30n w=0.17u
MM27 net166 net111 VDD VDD pch_mac l=30n w=0.17u
MM50 net111 mq VDD VDD pch_mac l=30n w=0.17u
MM29 net57 SI VDD VDD pch_mac l=30n w=100n
MM28 net54 net139 net57 VDD pch_mac l=30n w=100n
MM24 net58 SE VDD VDD pch_mac l=30n w=0.21u
MM23 net54 D net58 VDD pch_mac l=30n w=0.21u
MM22 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM19 net139 SE VDD VDD pch_mac l=30n w=0.21u
MM21 mq_x clkb net54 VDD pch_mac l=30n w=0.17u
MM20 clkb CPN VDD VDD pch_mac l=30n w=0.17u
MM60 net89 net166 VDD VDD pch_mac l=30n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM79 mq_x clkbb net89 VDD pch_mac l=30n w=0.17u
MM13 mq mq_x VDD VDD pch_mac l=30n w=0.17u
MM10 mq SDN VDD VDD pch_mac l=30n w=0.22u
MM4 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM4_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM8 net135 SDN VDD VDD pch_mac l=30n w=0.17u
MM30 net135 clkb qf VDD pch_mac l=30n w=0.17u
MM6 net135 qf_x VDD VDD pch_mac l=30n w=0.17u
MM2 QN net135 VDD VDD pch_mac l=30n w=0.17u 
MM2_2 QN net135 VDD VDD pch_mac l=30n w=0.17u 
MM33 net104 net111 VSS VSS nch_mac l=30n w=0.14u
MM31 qf clkb net104 VSS nch_mac l=30n w=0.22u
MM26 net166 net111 VSS VSS nch_mac l=30n w=0.14u
MM49 net111 mq VSS VSS nch_mac l=30n w=0.14u
MM15 net139 SE VSS VSS nch_mac l=30n w=0.22u
MM17 net143 SI VSS VSS nch_mac l=30n w=0.12u
MM16 net155 D net148 VSS nch_mac l=30n w=0.22u
MM0 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM18 net155 SE net143 VSS nch_mac l=30n w=0.12u
MM1 mq_x clkbb net155 VSS nch_mac l=30n w=0.14u
MM11 clkb CPN VSS VSS nch_mac l=30n w=0.14u
MM65 net172 net166 VSS VSS nch_mac l=30n w=0.14u
MM64 mq_x clkb net172 VSS nch_mac l=30n w=0.14u
MM76 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM12 net148 net139 VSS VSS nch_mac l=30n w=0.22u
MM5 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM5_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM3 QN net135 VSS VSS nch_mac l=30n w=0.14u 
MM3_2 QN net135 VSS VSS nch_mac l=30n w=0.14u 
MM9 net127 qf_x VSS VSS nch_mac l=30n w=0.14u
MM14 net184 mq_x VSS VSS nch_mac l=30n w=0.14u
MM25 mq SDN net184 VSS nch_mac l=30n w=0.14u
MM7 net135 SDN net127 VSS nch_mac l=30n w=0.14u
MM32 net135 clkbb qf VSS nch_mac l=30n w=0.22u
.ENDS
.SUBCKT SDFSYNCND2 SI D SE CP CDN Q QN VDD VSS
MM6 qf clkbb net0154 VSS nch_mac l=30n w=0.14u
MM7 net0154 net0232 VSS VSS nch_mac l=30n w=0.14u
MM12 net0171 SE net0172 VSS nch_mac l=30n w=0.12u
MM27 net0171 D net0187 VSS nch_mac l=30n w=0.22u
MM14 net0183 SE VSS VSS nch_mac l=30n w=0.22u
MM0 net0232 net0301 VSS VSS nch_mac l=30n w=0.14u
MM2 net0200 net0232 VSS VSS nch_mac l=30n w=0.14u
MM11 net0172 SI VSS VSS nch_mac l=30n w=0.12u
MM26 net0156 CDN net0148 VSS nch_mac l=30n w=0.14u
MM46 mq_x clkb net0171 VSS nch_mac l=30n w=0.14u
MM47 net0187 net0183 VSS VSS nch_mac l=30n w=0.22u
MM28 mq_x clkbb net0156 VSS nch_mac l=30n w=0.14u
MM73 net102 qf_x VSS VSS nch_mac l=30n w=0.14u
MM23 net102 clkb qf VSS nch_mac l=30n w=0.14u
MM69 QN net102 VSS VSS nch_mac l=30n w=0.14u 
MM69_2 QN net102 VSS VSS nch_mac l=30n w=0.14u 
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM29 net0148 net0200 VSS VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM76 qf_x qf net150 VSS nch_mac l=30n w=0.14u
MM49 net0301 mq_x VSS VSS nch_mac l=30n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM75 net150 CDN VSS VSS nch_mac l=30n w=0.14u
MM3 net0200 net0232 VDD VDD pch_mac l=30n w=0.17u
MM9 qf clkb net0236 VDD pch_mac l=30n w=0.17u
MM10 net0236 net0232 VDD VDD pch_mac l=30n w=0.17u
MM1 net0232 net0301 VDD VDD pch_mac l=30n w=0.17u
MM70 QN net102 VDD VDD pch_mac l=30n w=0.335u 
MM70_2 QN net102 VDD VDD pch_mac l=30n w=0.335u 
MM74 net102 qf_x VDD VDD pch_mac l=30n w=0.335u
MM5 net0234 CDN VDD VDD pch_mac l=30n w=0.17u
MM50 net0301 mq_x VDD VDD pch_mac l=30n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM13 net102 clkbb qf VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM16 net0183 SE VDD VDD pch_mac l=30n w=0.21u
MM45 mq_x clkbb net0262 VDD pch_mac l=30n w=0.17u
MM44 net0262 D net0266 VDD pch_mac l=30n w=0.21u
MM15 mq_x clkb net0234 VDD pch_mac l=30n w=0.17u
MM8 net0234 net0200 VDD VDD pch_mac l=30n w=0.17u
MM17 net0266 SE VDD VDD pch_mac l=30n w=0.21u
MM18 net0262 net0183 net0258 VDD pch_mac l=30n w=100n
MM19 net0258 SI VDD VDD pch_mac l=30n w=100n
.ENDS
.SUBCKT SDFSYNCNQD2 SI D SE CP CDN Q VDD VSS
MM19 net13 SI VDD VDD pch_mac l=30n w=0.12u
MM18 net17 net41 net13 VDD pch_mac l=30n w=0.12u
MM17 net21 SE VDD VDD pch_mac l=30n w=0.21u
MM8 net73 net113 VDD VDD pch_mac l=30n w=0.17u
MM15 mq_x clkb net73 VDD pch_mac l=30n w=0.17u
MM44 net17 D net21 VDD pch_mac l=30n w=0.21u
MM45 mq_x clkbb net17 VDD pch_mac l=30n w=0.17u
MM16 net41 SE VDD VDD pch_mac l=30n w=0.21u
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM13 net53 clkbb qf VDD pch_mac l=30n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM78 qf_x CDN VDD VDD pch_mac l=30n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM50 net69 mq_x VDD VDD pch_mac l=30n w=0.17u
MM5 net73 CDN VDD VDD pch_mac l=30n w=0.17u
MM74 net53 qf_x VDD VDD pch_mac l=30n w=0.335u
MM1 net154 net69 VDD VDD pch_mac l=30n w=0.17u
MM10 net81 net154 VDD VDD pch_mac l=30n w=0.17u
MM9 qf clkb net81 VDD pch_mac l=30n w=0.17u
MM3 net113 net154 VDD VDD pch_mac l=30n w=0.17u
MM75 net107 CDN VSS VSS nch_mac l=30n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM49 net69 mq_x VSS VSS nch_mac l=30n w=0.14u
MM76 qf_x qf net107 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM29 net114 net113 VSS VSS nch_mac l=30n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM23 net122 clkb qf VSS nch_mac l=30n w=0.14u
MM73 net122 qf_x VSS VSS nch_mac l=30n w=0.14u
MM28 mq_x clkbb net131 VSS nch_mac l=30n w=0.14u
MM47 net134 net41 VSS VSS nch_mac l=30n w=0.22u
MM46 mq_x clkb net166 VSS nch_mac l=30n w=0.14u
MM26 net131 CDN net114 VSS nch_mac l=30n w=0.14u
MM11 net167 SI VSS VSS nch_mac l=30n w=0.12u
MM2 net113 net154 VSS VSS nch_mac l=30n w=0.14u
MM0 net154 net69 VSS VSS nch_mac l=30n w=0.14u
MM14 net41 SE VSS VSS nch_mac l=30n w=0.22u
MM27 net166 D net134 VSS nch_mac l=30n w=0.22u
MM12 net166 SE net167 VSS nch_mac l=30n w=0.12u
MM7 net175 net154 VSS VSS nch_mac l=30n w=0.14u
MM6 qf clkbb net175 VSS nch_mac l=30n w=0.14u
.ENDS
.SUBCKT SDFSYNCSND2 SI D SE CP CDN SDN Q QN VDD VSS
MM21 net18 net23 VDD VDD pch_mac l=30n w=0.17u
MM16 net167 net23 VDD VDD pch_mac l=30n w=0.17u
MM15 net23 mq VDD VDD pch_mac l=30n w=0.17u
MM20 qf clkb net18 VDD pch_mac l=30n w=0.17u
MM1 mq net59 VDD VDD pch_mac l=30n w=0.17u
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM43 net90 SE VDD VDD pch_mac l=30n w=0.21u
MM11 net91 CDN VDD VDD pch_mac l=30n w=0.17u
MM14 net132 clkbb qf VDD pch_mac l=30n w=0.17u
MM44 net55 D net90 VDD pch_mac l=30n w=0.21u
MM77 qf_x CDN VDD VDD pch_mac l=30n w=0.33u
MM78 qf_x qf VDD VDD pch_mac l=30n w=0.33u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM12 net59 clkb net91 VDD pch_mac l=30n w=0.17u
MM0 mq SDN VDD VDD pch_mac l=30n w=0.17u
MM41 net58 SI VDD VDD pch_mac l=30n w=100n
MM13 net91 net167 VDD VDD pch_mac l=30n w=0.17u
MM58 net172 SE VDD VDD pch_mac l=30n w=0.21u
MM70 QN net132 VDD VDD pch_mac l=30n w=0.17u 
MM70_2 QN net132 VDD VDD pch_mac l=30n w=0.17u 
MM45 net59 clkbb net55 VDD pch_mac l=30n w=0.17u
MM42 net55 net172 net58 VDD pch_mac l=30n w=100n
MM4 net132 qf_x VDD VDD pch_mac l=30n w=0.33u
MM5 net132 SDN VDD VDD pch_mac l=30n w=0.33u
MM18 qf clkbb net108 VSS nch_mac l=30n w=0.14u
MM49 net23 mq VSS VSS nch_mac l=30n w=0.14u
MM17 net167 net23 VSS VSS nch_mac l=30n w=0.14u
MM19 net108 net23 VSS VSS nch_mac l=30n w=0.14u
MM75 net145 qf VSS VSS nch_mac l=30n w=0.275u
MM47 net160 D net164 VSS nch_mac l=30n w=0.22u
MM51 net161 SI VSS VSS nch_mac l=30n w=0.12u
MM46 net59 clkb net160 VSS nch_mac l=30n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM76 qf_x CDN net145 VSS nch_mac l=30n w=0.275u
MM9 net59 clkbb net177 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM8 net177 CDN net181 VSS nch_mac l=30n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM57 net172 SE VSS VSS nch_mac l=30n w=0.22u
MM10 net181 net167 VSS VSS nch_mac l=30n w=0.14u
MM48 net164 net172 VSS VSS nch_mac l=30n w=0.22u
MM69 QN net132 VSS VSS nch_mac l=30n w=0.14u 
MM69_2 QN net132 VSS VSS nch_mac l=30n w=0.14u 
MM50 net132 clkb qf VSS nch_mac l=30n w=0.14u
MM2 mq SDN net157 VSS nch_mac l=30n w=0.14u
MM52 net160 SE net161 VSS nch_mac l=30n w=0.12u
MM6 net132 SDN net125 VSS nch_mac l=30n w=0.275u
MM3 net157 net59 VSS VSS nch_mac l=30n w=0.14u
MM7 net125 qf_x VSS VSS nch_mac l=30n w=0.275u
.ENDS
.SUBCKT SDFSYNCSNQD2 SI D SE CP CDN SDN Q VDD VSS
MM7 net11 qf_x VSS VSS nch_mac l=30n w=0.14u
MM3 net15 net71 VSS VSS nch_mac l=30n w=0.14u
MM6 net0182 SDN net11 VSS nch_mac l=30n w=0.14u
MM52 net23 SE net24 VSS nch_mac l=30n w=0.12u
MM2 mq SDN net15 VSS nch_mac l=30n w=0.14u
MM50 net0182 clkb qf VSS nch_mac l=30n w=0.14u
MM48 net35 net43 VSS VSS nch_mac l=30n w=0.22u
MM10 net39 net38 VSS VSS nch_mac l=30n w=0.14u
MM57 net43 SE VSS VSS nch_mac l=30n w=0.22u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM8 net51 CDN net39 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM9 net71 clkbb net51 VSS nch_mac l=30n w=0.14u
MM76 qf_x qf net83 VSS nch_mac l=30n w=0.14u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM46 net71 clkb net23 VSS nch_mac l=30n w=0.14u
MM51 net24 SI VSS VSS nch_mac l=30n w=0.12u
MM47 net23 D net35 VSS nch_mac l=30n w=0.22u
MM75 net83 CDN VSS VSS nch_mac l=30n w=0.14u
MM19 net100 net182 VSS VSS nch_mac l=30n w=0.14u
MM17 net38 net182 VSS VSS nch_mac l=30n w=0.14u
MM49 net182 mq VSS VSS nch_mac l=30n w=0.14u
MM18 qf clkbb net100 VSS nch_mac l=30n w=0.14u
MM5 net31 SDN VDD VDD pch_mac l=30n w=0.335u
MM4 net31 qf_x VDD VDD pch_mac l=30n w=0.335u
MM42 net110 net43 net126 VDD pch_mac l=30n w=0.12u
MM45 net71 clkbb net110 VDD pch_mac l=30n w=0.17u
MM58 net43 SE VDD VDD pch_mac l=30n w=0.21u
MM13 net158 net38 VDD VDD pch_mac l=30n w=0.17u
MM41 net126 SI VDD VDD pch_mac l=30n w=0.12u
MM0 mq SDN VDD VDD pch_mac l=30n w=0.17u
MM12 net71 clkb net158 VDD pch_mac l=30n w=0.17u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM78 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM77 qf_x CDN VDD VDD pch_mac l=30n w=0.17u
MM44 net110 D net153 VDD pch_mac l=30n w=0.21u
MM14 net31 clkbb qf VDD pch_mac l=30n w=0.17u
MM11 net158 CDN VDD VDD pch_mac l=30n w=0.17u
MM43 net153 SE VDD VDD pch_mac l=30n w=0.21u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM1 mq net71 VDD VDD pch_mac l=30n w=0.17u
MM20 qf clkb net181 VDD pch_mac l=30n w=0.17u
MM15 net182 mq VDD VDD pch_mac l=30n w=0.17u
MM16 net38 net182 VDD VDD pch_mac l=30n w=0.17u
MM21 net181 net182 VDD VDD pch_mac l=30n w=0.17u
.ENDS
.SUBCKT SDFSYND2 SI D SE CP Q QN VDD VSS
MM0 net0240 net0176 VSS VSS nch_mac l=30n w=0.14u
MM5 net0188 net0240 VSS VSS nch_mac l=30n w=0.14u
MM47 net61 D net0177 VSS nch_mac l=30n w=0.22u
MM51 net13 SI VSS VSS nch_mac l=30n w=0.12u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM49 net0176 mq_x VSS VSS nch_mac l=30n w=0.14u
MM46 mq_x clkb net61 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM26 net0136 net0188 VSS VSS nch_mac l=30n w=0.14u
MM57 net0241 SE VSS VSS nch_mac l=30n w=0.22u
MM28 mq_x clkbb net0136 VSS nch_mac l=30n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM30 net49 clkb qf VSS nch_mac l=30n w=0.14u
MM48 net0177 net0241 VSS VSS nch_mac l=30n w=0.22u
MM7 net0157 net0240 VSS VSS nch_mac l=30n w=0.14u
MM52 net61 SE net13 VSS nch_mac l=30n w=0.12u
MM2 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM69 QN net49 VSS VSS nch_mac l=30n w=0.14u 
MM69_2 QN net49 VSS VSS nch_mac l=30n w=0.14u 
MM73 net49 qf_x VSS VSS nch_mac l=30n w=0.14u
MM9 qf clkbb net0157 VSS nch_mac l=30n w=0.14u
MM4 net0188 net0240 VDD VDD pch_mac l=30n w=0.17u
MM12 net0236 net0240 VDD VDD pch_mac l=30n w=0.17u
MM13 qf clkb net0236 VDD pch_mac l=30n w=0.17u
MM3 net0240 net0176 VDD VDD pch_mac l=30n w=0.17u
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM43 net53 SE VDD VDD pch_mac l=30n w=0.21u
MM6 net0202 net0188 VDD VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM8 net49 clkbb qf VDD pch_mac l=30n w=0.17u
MM44 net125 D net53 VDD pch_mac l=30n w=0.21u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM50 net0176 mq_x VDD VDD pch_mac l=30n w=0.17u
MM41 net128 SI VDD VDD pch_mac l=30n w=0.12u
MM58 net0241 SE VDD VDD pch_mac l=30n w=0.21u
MM45 mq_x clkbb net125 VDD pch_mac l=30n w=0.17u
MM42 net125 net0241 net128 VDD pch_mac l=30n w=0.12u
MM16 mq_x clkb net0202 VDD pch_mac l=30n w=0.17u
MM1 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM74 net49 qf_x VDD VDD pch_mac l=30n w=0.17u
MM70 QN net49 VDD VDD pch_mac l=30n w=0.17u 
MM70_2 QN net49 VDD VDD pch_mac l=30n w=0.17u 
.ENDS
.SUBCKT SDFSYNQD2 SI D SE CP Q VDD VSS
MM0 net0240 net0176 VSS VSS nch_mac l=30n w=0.14u
MM5 net0188 net0240 VSS VSS nch_mac l=30n w=0.14u
MM47 net61 D net0177 VSS nch_mac l=30n w=0.22u
MM51 net13 SI VSS VSS nch_mac l=30n w=0.12u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM49 net0176 mq_x VSS VSS nch_mac l=30n w=0.14u
MM46 mq_x clkb net61 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM26 net0136 net0188 VSS VSS nch_mac l=30n w=0.14u
MM57 net0241 SE VSS VSS nch_mac l=30n w=0.22u
MM28 mq_x clkbb net0136 VSS nch_mac l=30n w=0.14u
MM71 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM71_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM30 net49 clkb qf VSS nch_mac l=30n w=0.14u
MM48 net0177 net0241 VSS VSS nch_mac l=30n w=0.22u
MM7 net0157 net0240 VSS VSS nch_mac l=30n w=0.14u
MM52 net61 SE net13 VSS nch_mac l=30n w=0.12u
MM2 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM73 net49 qf_x VSS VSS nch_mac l=30n w=0.14u
MM9 qf clkbb net0157 VSS nch_mac l=30n w=0.14u
MM4 net0188 net0240 VDD VDD pch_mac l=30n w=0.17u
MM12 net0236 net0240 VDD VDD pch_mac l=30n w=0.17u
MM13 qf clkb net0236 VDD pch_mac l=30n w=0.17u
MM3 net0240 net0176 VDD VDD pch_mac l=30n w=0.17u
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM43 net53 SE VDD VDD pch_mac l=30n w=0.21u
MM6 net0202 net0188 VDD VDD pch_mac l=30n w=0.17u
MM72 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM72_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM8 net0421 clkbb qf VDD pch_mac l=30n w=0.17u
MM44 net125 D net53 VDD pch_mac l=30n w=0.21u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM50 net0176 mq_x VDD VDD pch_mac l=30n w=0.17u
MM41 net128 SI VDD VDD pch_mac l=30n w=0.12u
MM58 net0241 SE VDD VDD pch_mac l=30n w=0.21u
MM45 mq_x clkbb net125 VDD pch_mac l=30n w=0.17u
MM42 net125 net0241 net128 VDD pch_mac l=30n w=0.12u
MM16 mq_x clkb net0202 VDD pch_mac l=30n w=0.17u
MM1 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM74 net0421 qf_x VDD VDD pch_mac l=30n w=0.17u
.ENDS
.SUBCKT SDFSYNQND2 SI D SE CP QN VDD VSS
MM0 net0240 net0176 VSS VSS nch_mac l=30n w=0.14u
MM5 net0188 net0240 VSS VSS nch_mac l=30n w=0.14u
MM47 net61 D net0177 VSS nch_mac l=30n w=0.22u
MM51 net13 SI VSS VSS nch_mac l=30n w=0.12u
MM53 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM49 net0176 mq_x VSS VSS nch_mac l=30n w=0.14u
MM46 mq_x clkb net61 VSS nch_mac l=30n w=0.14u
MM55 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM26 net0136 net0188 VSS VSS nch_mac l=30n w=0.14u
MM57 net0241 SE VSS VSS nch_mac l=30n w=0.22u
MM28 mq_x clkbb net0136 VSS nch_mac l=30n w=0.14u
MM71 QN qf VSS VSS nch_mac l=30n w=0.14u 
MM71_2 QN qf VSS VSS nch_mac l=30n w=0.14u 
MM30 net49 clkb qf VSS nch_mac l=30n w=0.14u
MM48 net0177 net0241 VSS VSS nch_mac l=30n w=0.22u
MM7 net0157 net0240 VSS VSS nch_mac l=30n w=0.14u
MM52 net61 SE net13 VSS nch_mac l=30n w=0.12u
MM2 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM73 net49 qf_x VSS VSS nch_mac l=30n w=0.14u
MM9 qf clkbb net0157 VSS nch_mac l=30n w=0.14u
MM4 net0188 net0240 VDD VDD pch_mac l=30n w=0.17u
MM12 net0236 net0240 VDD VDD pch_mac l=30n w=0.17u
MM13 qf clkb net0236 VDD pch_mac l=30n w=0.17u
MM3 net0240 net0176 VDD VDD pch_mac l=30n w=0.17u
MM54 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM43 net53 SE VDD VDD pch_mac l=30n w=0.21u
MM6 net0202 net0188 VDD VDD pch_mac l=30n w=0.17u
MM72 QN qf VDD VDD pch_mac l=30n w=0.17u 
MM72_2 QN qf VDD VDD pch_mac l=30n w=0.17u 
MM8 net0253 clkbb qf VDD pch_mac l=30n w=0.17u
MM44 net125 D net53 VDD pch_mac l=30n w=0.21u
MM56 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM50 net0176 mq_x VDD VDD pch_mac l=30n w=0.17u
MM41 net128 SI VDD VDD pch_mac l=30n w=0.12u
MM58 net0241 SE VDD VDD pch_mac l=30n w=0.21u
MM45 mq_x clkbb net125 VDD pch_mac l=30n w=0.17u
MM42 net125 net0241 net128 VDD pch_mac l=30n w=0.12u
MM16 mq_x clkb net0202 VDD pch_mac l=30n w=0.17u
MM1 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM74 net0253 qf_x VDD VDD pch_mac l=30n w=0.17u
.ENDS
.SUBCKT SDFSYNSND2 SI D SE CP SDN Q QN VDD VSS
MM35 net10 net111 VDD VDD pch_mac l=30n w=0.17u
MM34 qf clkb net10 VDD pch_mac l=30n w=0.17u
MM27 net166 net111 VDD VDD pch_mac l=30n w=0.17u
MM50 net111 mq VDD VDD pch_mac l=30n w=0.17u
MM29 net57 SI VDD VDD pch_mac l=30n w=0.12u
MM28 net54 net139 net57 VDD pch_mac l=30n w=0.12u
MM24 net58 SE VDD VDD pch_mac l=30n w=0.21u
MM23 net54 D net58 VDD pch_mac l=30n w=0.21u
MM22 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM19 net139 SE VDD VDD pch_mac l=30n w=0.21u
MM21 mq_x clkbb net54 VDD pch_mac l=30n w=0.17u
MM20 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM60 net89 net166 VDD VDD pch_mac l=30n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM79 mq_x clkb net89 VDD pch_mac l=30n w=0.17u
MM13 mq mq_x VDD VDD pch_mac l=30n w=0.17u
MM10 mq SDN VDD VDD pch_mac l=30n w=0.22u
MM4 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM4_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM8 net135 SDN VDD VDD pch_mac l=30n w=0.17u
MM30 net135 clkbb qf VDD pch_mac l=30n w=0.17u
MM6 net135 qf_x VDD VDD pch_mac l=30n w=0.17u
MM2 QN net135 VDD VDD pch_mac l=30n w=0.17u 
MM2_2 QN net135 VDD VDD pch_mac l=30n w=0.17u 
MM33 net104 net111 VSS VSS nch_mac l=30n w=0.14u
MM31 qf clkbb net104 VSS nch_mac l=30n w=0.22u
MM26 net166 net111 VSS VSS nch_mac l=30n w=0.14u
MM49 net111 mq VSS VSS nch_mac l=30n w=0.14u
MM15 net139 SE VSS VSS nch_mac l=30n w=0.22u
MM17 net143 SI VSS VSS nch_mac l=30n w=0.12u
MM16 net155 D net148 VSS nch_mac l=30n w=0.22u
MM0 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM18 net155 SE net143 VSS nch_mac l=30n w=0.12u
MM1 mq_x clkb net155 VSS nch_mac l=30n w=0.14u
MM11 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM65 net172 net166 VSS VSS nch_mac l=30n w=0.14u
MM64 mq_x clkbb net172 VSS nch_mac l=30n w=0.14u
MM76 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM12 net148 net139 VSS VSS nch_mac l=30n w=0.22u
MM5 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM5_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM3 QN net135 VSS VSS nch_mac l=30n w=0.14u 
MM3_2 QN net135 VSS VSS nch_mac l=30n w=0.14u 
MM9 net127 qf_x VSS VSS nch_mac l=30n w=0.14u
MM14 net184 mq_x VSS VSS nch_mac l=30n w=0.14u
MM25 mq SDN net184 VSS nch_mac l=30n w=0.14u
MM7 net135 SDN net127 VSS nch_mac l=30n w=0.14u
MM32 net135 clkb qf VSS nch_mac l=30n w=0.22u
.ENDS
.SUBCKT SDFSYNSNQD2 SI D SE CP SDN Q VDD VSS
MM35 net10 net111 VDD VDD pch_mac l=30n w=0.17u
MM34 qf clkb net10 VDD pch_mac l=30n w=0.17u
MM27 net166 net111 VDD VDD pch_mac l=30n w=0.17u
MM50 net111 mq VDD VDD pch_mac l=30n w=0.17u
MM29 net57 SI VDD VDD pch_mac l=30n w=100n
MM28 net54 net139 net57 VDD pch_mac l=30n w=100n
MM24 net58 SE VDD VDD pch_mac l=30n w=0.21u
MM23 net54 D net58 VDD pch_mac l=30n w=0.21u
MM22 clkbb clkb VDD VDD pch_mac l=30n w=0.17u
MM19 net139 SE VDD VDD pch_mac l=30n w=0.21u
MM21 mq_x clkbb net54 VDD pch_mac l=30n w=0.17u
MM20 clkb CP VDD VDD pch_mac l=30n w=0.17u
MM60 net89 net166 VDD VDD pch_mac l=30n w=0.17u
MM77 qf_x qf VDD VDD pch_mac l=30n w=0.17u
MM79 mq_x clkb net89 VDD pch_mac l=30n w=0.17u
MM13 mq mq_x VDD VDD pch_mac l=30n w=0.17u
MM10 mq SDN VDD VDD pch_mac l=30n w=0.22u
MM4 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM4_2 Q qf_x VDD VDD pch_mac l=30n w=0.17u 
MM8 net135 SDN VDD VDD pch_mac l=30n w=0.17u
MM30 net135 clkbb qf VDD pch_mac l=30n w=0.17u
MM6 net135 qf_x VDD VDD pch_mac l=30n w=0.17u
MM33 net104 net111 VSS VSS nch_mac l=30n w=0.14u
MM31 qf clkbb net104 VSS nch_mac l=30n w=0.22u
MM26 net166 net111 VSS VSS nch_mac l=30n w=0.14u
MM49 net111 mq VSS VSS nch_mac l=30n w=0.14u
MM15 net139 SE VSS VSS nch_mac l=30n w=0.22u
MM17 net143 SI VSS VSS nch_mac l=30n w=0.12u
MM16 net155 D net148 VSS nch_mac l=30n w=0.22u
MM0 clkbb clkb VSS VSS nch_mac l=30n w=0.14u
MM18 net155 SE net143 VSS nch_mac l=30n w=0.12u
MM1 mq_x clkb net155 VSS nch_mac l=30n w=0.14u
MM11 clkb CP VSS VSS nch_mac l=30n w=0.14u
MM65 net172 net166 VSS VSS nch_mac l=30n w=0.14u
MM64 mq_x clkbb net172 VSS nch_mac l=30n w=0.14u
MM76 qf_x qf VSS VSS nch_mac l=30n w=0.14u
MM12 net148 net139 VSS VSS nch_mac l=30n w=0.22u
MM5 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM5_2 Q qf_x VSS VSS nch_mac l=30n w=0.14u 
MM9 net127 qf_x VSS VSS nch_mac l=30n w=0.14u
MM14 net184 mq_x VSS VSS nch_mac l=30n w=0.14u
MM25 mq SDN net184 VSS nch_mac l=30n w=0.14u
MM7 net135 SDN net127 VSS nch_mac l=30n w=0.14u
MM32 net135 clkb qf VSS nch_mac l=30n w=0.22u
.ENDS
.SUBCKT GAN2MCOD2 A1 A2 Z VDD VSS
MM9 net14 A2 VSS VSS nch_mac l=0.03u w=0.14u
MM8 net26 A1 net14 VSS nch_mac l=0.03u w=0.14u
MM5 Z net26 VSS VSS nch_mac l=0.03u w=0.14u 
MM5_2 Z net26 VSS VSS nch_mac l=0.03u w=0.14u 
MM6 net26 A1 VDD VDD pch_mac l=0.03u w=0.17u
MM7 net26 A2 VDD VDD pch_mac l=0.03u w=0.17u
MM4 Z net26 VDD VDD pch_mac l=0.03u w=0.17u 
MM4_2 Z net26 VDD VDD pch_mac l=0.03u w=0.17u 
.ENDS
.SUBCKT GAOI21MCOD2 A1 A2 B ZN VDD VSS
MM9 VSS B VSS VSS nch_mac l=0.03u w=0.14u
MM5 ZN A1 net027 VSS nch_mac l=0.03u w=0.14u
MM4 net027 A2 VSS VSS nch_mac l=0.03u w=0.14u
MM2 net7 A2 VSS VSS nch_mac l=0.03u w=0.14u
MM1 ZN A1 net7 VSS nch_mac l=0.03u w=0.14u
MM0 ZN B VSS VSS nch_mac l=0.03u w=0.14u
MM8 VDD B VDD VDD pch_mac l=0.03u w=0.17u
MM7 net30 B VDD VDD pch_mac l=0.03u w=0.17u
MM6 ZN A2 net30 VDD pch_mac l=0.03u w=0.17u 
MM6_2 ZN A2 net30 VDD pch_mac l=0.03u w=0.17u 
MM3 ZN A1 net30 VDD pch_mac l=0.03u w=0.17u 
MM3_2 ZN A1 net30 VDD pch_mac l=0.03u w=0.17u 
.ENDS
.SUBCKT GBUFFMCOD2 I Z VDD VSS
MM26 VSS I VSS VSS nch_mac l=0.03u w=0.14u
MM0 Z net9 VSS VSS nch_mac l=0.03u w=0.14u 
MM0_2 Z net9 VSS VSS nch_mac l=0.03u w=0.14u 
MM5 net9 I VSS VSS nch_mac l=0.03u w=0.14u
MM24 VDD I VDD VDD pch_mac l=0.03u w=0.17u
MM1 Z net9 VDD VDD pch_mac l=0.03u w=0.17u 
MM1_2 Z net9 VDD VDD pch_mac l=0.03u w=0.17u 
MM4 net9 I VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GINVMCOD2 I ZN VDD VSS
MM0 ZN I VDD VDD pch_mac l=0.03u w=0.17u 
MM0_2 ZN I VDD VDD pch_mac l=0.03u w=0.17u 
MM6 net37 net37 net37 VDD pch_mac l=0.03u w=0.17u
MM5 net37 net35 net37 VDD pch_mac l=0.03u w=0.17u
MM4 net35 net35 net35 VSS nch_mac l=0.03u w=0.14u
MM1 ZN I VSS VSS nch_mac l=0.03u w=0.14u 
MM1_2 ZN I VSS VSS nch_mac l=0.03u w=0.14u 
MM8 net35 net37 net35 VSS nch_mac l=0.03u w=0.14u
.ENDS
.SUBCKT GMUX2MCOD2 I0 I1 S Z VDD VSS
MM19 VSS S VSS VSS nch_mac l=0.03u w=0.14u
MM6 nn1 I1 VSS VSS nch_mac l=0.03u w=0.14u
MM18 VSS I0 VSS VSS nch_mac l=0.03u w=0.14u
MM9 sb S VSS VSS nch_mac l=0.03u w=0.14u
MM2 net62 I0 VSS VSS nch_mac l=0.03u w=0.14u
MM7 net53 S nn1 VSS nch_mac l=0.03u w=0.14u
MM12 Z net53 VSS VSS nch_mac l=0.03u w=0.14u 
MM12_2 Z net53 VSS VSS nch_mac l=0.03u w=0.14u 
MM0 net53 sb net62 VSS nch_mac l=0.03u w=0.14u
MM16 nn1 sb nn1 VSS nch_mac l=0.03u w=0.14u
MM10 VDD I0 VDD VDD pch_mac l=0.03u w=0.17u
MM17 pp1 sb pp1 VDD pch_mac l=0.03u w=0.17u
MM11 VDD S VDD VDD pch_mac l=0.03u w=0.17u
MM14 net93 I1 VDD VDD pch_mac l=0.03u w=0.17u
MM8 sb S VDD VDD pch_mac l=0.03u w=0.17u
MM13 Z net53 VDD VDD pch_mac l=0.03u w=0.17u 
MM13_2 Z net53 VDD VDD pch_mac l=0.03u w=0.17u 
MM1 net53 S pp1 VDD pch_mac l=0.03u w=0.17u
MM3 pp1 I0 VDD VDD pch_mac l=0.03u w=0.17u
MM5 net53 sb net93 VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GMUX2NMCOD2 I0 I1 S ZN VDD VSS
MM6 net0148 I1 VSS VSS nch_mac l=0.03u w=0.14u
MM17 VSS S VSS VSS nch_mac l=0.03u w=0.14u
MM19 n1 S n1 VSS nch_mac l=0.03u w=0.14u
MM12 ZN net88 VSS VSS nch_mac l=0.03u w=0.14u 
MM12_2 ZN net88 VSS VSS nch_mac l=0.03u w=0.14u 
MM9 sn S VSS VSS nch_mac l=0.03u w=0.14u
MM7 zb S net0148 VSS nch_mac l=0.03u w=0.14u
MM2 n1 I0 VSS VSS nch_mac l=0.03u w=0.14u
MM0 zb sn n1 VSS nch_mac l=0.03u w=0.14u
MM11 net88 zb VSS VSS nch_mac l=0.03u w=0.14u
MM13 ZN net88 VDD VDD pch_mac l=0.03u w=0.17u 
MM13_2 ZN net88 VDD VDD pch_mac l=0.03u w=0.17u 
MM1 zb S net0190 VDD pch_mac l=0.03u w=0.17u
MM5 zb sn pp1 VDD pch_mac l=0.03u w=0.17u
MM8 sn S VDD VDD pch_mac l=0.03u w=0.17u
MM3 net0190 I0 VDD VDD pch_mac l=0.03u w=0.17u
MM10 net88 zb VDD VDD pch_mac l=0.03u w=0.17u
MM18 pp1 S pp1 VDD pch_mac l=0.03u w=0.17u
MM16 VDD S VDD VDD pch_mac l=0.03u w=0.17u
MM4 pp1 I1 VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GND2MCOD2 A1 A2 ZN VDD VSS
MM0 net33 A2 VSS VSS nch_mac l=0.03u w=0.14u
MM3 ZN A1 net33 VSS nch_mac l=0.03u w=0.14u
MM4 VSS A2 VSS VSS nch_mac l=0.03u w=0.14u 
MM4_2 VSS A2 VSS VSS nch_mac l=0.03u w=0.14u 
MM7 net28 A2 VSS VSS nch_mac l=0.03u w=0.14u
MM6 ZN A1 net28 VSS nch_mac l=0.03u w=0.14u
MM5 VDD A2 VDD VDD pch_mac l=0.03u w=0.17u 
MM5_2 VDD A2 VDD VDD pch_mac l=0.03u w=0.17u 
MM2 ZN A1 VDD VDD pch_mac l=0.03u w=0.17u 
MM2_2 ZN A1 VDD VDD pch_mac l=0.03u w=0.17u 
MM1 ZN A2 VDD VDD pch_mac l=0.03u w=0.17u 
MM1_2 ZN A2 VDD VDD pch_mac l=0.03u w=0.17u 
.ENDS
.SUBCKT GND3MCOD2 A1 A2 A3 ZN VDD VSS
MM7 net33 A2 net61 VSS nch_mac l=0.03u w=0.14u
MM8 ZN A3 net33 VSS nch_mac l=0.03u w=0.14u
MM2 net41 A1 VSS VSS nch_mac l=0.03u w=0.14u
MM1 net46 A2 net41 VSS nch_mac l=0.03u w=0.14u
MM0 ZN A3 net46 VSS nch_mac l=0.03u w=0.14u
MM6 net61 A1 VSS VSS nch_mac l=0.03u w=0.14u
MM4 ZN A1 VDD VDD pch_mac l=0.03u w=0.17u 
MM4_2 ZN A1 VDD VDD pch_mac l=0.03u w=0.17u 
MM5 ZN A3 VDD VDD pch_mac l=0.03u w=0.17u 
MM5_2 ZN A3 VDD VDD pch_mac l=0.03u w=0.17u 
MM3 ZN A2 VDD VDD pch_mac l=0.03u w=0.17u 
MM3_2 ZN A2 VDD VDD pch_mac l=0.03u w=0.17u 
.ENDS
.SUBCKT GNR2MCOD2 A1 A2 ZN VDD VSS
MM1 ZN A1 VSS VSS nch_mac l=0.03u w=0.14u 
MM1_2 ZN A1 VSS VSS nch_mac l=0.03u w=0.14u 
MM0 ZN A2 VSS VSS nch_mac l=0.03u w=0.14u 
MM0_2 ZN A2 VSS VSS nch_mac l=0.03u w=0.14u 
MM3 ZN A2 net45 VDD pch_mac l=0.03u w=0.17u
MM6 net37 A1 VDD VDD pch_mac l=0.03u w=0.17u
MM4 ZN A2 net37 VDD pch_mac l=0.03u w=0.17u
MM2 net45 A1 VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GNR3MCOD2 A1 A2 A3 ZN VDD VSS
MM0 ZN A2 VSS VSS nch_mac l=0.03u w=0.14u 
MM0_2 ZN A2 VSS VSS nch_mac l=0.03u w=0.14u 
MM3 ZN A1 VSS VSS nch_mac l=0.03u w=0.14u 
MM3_2 ZN A1 VSS VSS nch_mac l=0.03u w=0.14u 
MM1 ZN A3 VSS VSS nch_mac l=0.03u w=0.14u 
MM1_2 ZN A3 VSS VSS nch_mac l=0.03u w=0.14u 
MM6 net56 A2 net44 VDD pch_mac l=0.03u w=0.17u 
MM6_2 net56 A2 net44 VDD pch_mac l=0.03u w=0.17u 
MM4 ZN A1 net56 VDD pch_mac l=0.03u w=0.17u 
MM4_2 ZN A1 net56 VDD pch_mac l=0.03u w=0.17u 
MM2 net44 A3 VDD VDD pch_mac l=0.03u w=0.17u 
MM2_2 net44 A3 VDD VDD pch_mac l=0.03u w=0.17u 
.ENDS
.SUBCKT GOAI21MCOD2 A1 A2 B ZN VDD VSS
MM8 net041 net041 net041 VSS nch_mac l=0.03u w=0.14u
MM9 net041 net035 net041 VSS nch_mac l=0.03u w=0.14u
MM3 net30 B VSS VSS nch_mac l=0.03u w=0.14u 
MM3_2 net30 B VSS VSS nch_mac l=0.03u w=0.14u 
MM58 ZN A2 net30 VSS nch_mac l=0.03u w=0.14u 
MM58_2 ZN A2 net30 VSS nch_mac l=0.03u w=0.14u 
MM2 ZN A1 net30 VSS nch_mac l=0.03u w=0.14u 
MM2_2 ZN A1 net30 VSS nch_mac l=0.03u w=0.14u 
MM6 net035 net041 net035 VDD pch_mac l=0.03u w=0.17u
MM7 net035 net035 net035 VDD pch_mac l=0.03u w=0.17u
MM4 ZN A1 net031 VDD pch_mac l=0.03u w=0.17u
MM5 net031 A2 VDD VDD pch_mac l=0.03u w=0.17u
MM59 ZN B VDD VDD pch_mac l=0.03u w=0.17u 
MM59_2 ZN B VDD VDD pch_mac l=0.03u w=0.17u 
MM0 ZN A1 net14 VDD pch_mac l=0.03u w=0.17u
MM1 net14 A2 VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GOR2MCOD2 A1 A2 Z VDD VSS
MM0 Z net26 VSS VSS nch_mac l=0.03u w=0.14u 
MM0_2 Z net26 VSS VSS nch_mac l=0.03u w=0.14u 
MM8 net26 A2 VSS VSS nch_mac l=0.03u w=0.14u
MM9 net26 A1 VSS VSS nch_mac l=0.03u w=0.14u
MM1 Z net26 VDD VDD pch_mac l=0.03u w=0.17u 
MM1_2 Z net26 VDD VDD pch_mac l=0.03u w=0.17u 
MM3 net26 A1 net13 VDD pch_mac l=0.03u w=0.17u
MM7 net13 A2 VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GXNR2MCOD2 A1 A2 ZN VDD VSS
MM12 a2n a1n a2n VSS nch_mac l=0.03u w=0.14u
MM11 net049 net051 net049 VSS nch_mac l=0.03u w=0.14u
MM10 net049 net049 net049 VSS nch_mac l=0.03u w=0.14u
MM3 net37 a1n net49 VSS nch_mac l=0.03u w=0.14u
MM1 net49 a2n VSS VSS nch_mac l=0.03u w=0.14u
MM6 ZN net37 VSS VSS nch_mac l=0.03u w=0.14u 
MM6_2 ZN net37 VSS VSS nch_mac l=0.03u w=0.14u 
MM0 a2n A2 VSS VSS nch_mac l=0.03u w=0.14u
MM17 a2n A1 net37 VSS nch_mac l=0.03u w=0.14u
MM8 a1n A1 VSS VSS nch_mac l=0.03u w=0.14u
MM13 pp1 a1n pp1 VDD pch_mac l=0.03u w=0.17u
MM4 net051 net051 net051 VDD pch_mac l=0.03u w=0.17u
MM5 net051 net049 net051 VDD pch_mac l=0.03u w=0.17u
MM15 net37 A1 pp1 VDD pch_mac l=0.03u w=0.17u
MM14 pp1 a2n VDD VDD pch_mac l=0.03u w=0.17u
MM7 ZN net37 VDD VDD pch_mac l=0.03u w=0.17u 
MM7_2 ZN net37 VDD VDD pch_mac l=0.03u w=0.17u 
MM2 a2n A2 VDD VDD pch_mac l=0.03u w=0.17u
MM16 a2n a1n net37 VDD pch_mac l=0.03u w=0.17u
MM9 a1n A1 VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT GXOR2MCOD2 A1 A2 Z VDD VSS
MM10 net054 net054 net054 VSS nch_mac l=0.03u w=0.14u
MM11 net054 net048 net054 VSS nch_mac l=0.03u w=0.14u
MM1 nn1 a2n VSS VSS nch_mac l=0.03u w=0.14u
MM3 zb A1 nn1 VSS nch_mac l=0.03u w=0.14u
MM8 a1n A1 VSS VSS nch_mac l=0.03u w=0.14u
MM0 a2n A2 VSS VSS nch_mac l=0.03u w=0.14u
MM6 Z zb VSS VSS nch_mac l=0.03u w=0.14u 
MM6_2 Z zb VSS VSS nch_mac l=0.03u w=0.14u 
MM17 zb a1n a2n VSS nch_mac l=0.03u w=0.14u
MM12 nn1 a1n nn1 VSS nch_mac l=0.03u w=0.14u
MM5 net048 net054 net048 VDD pch_mac l=0.03u w=0.17u
MM4 net048 net048 net048 VDD pch_mac l=0.03u w=0.17u
MM2 a2n A2 VDD VDD pch_mac l=0.03u w=0.17u
MM16 zb A1 a2n VDD pch_mac l=0.03u w=0.17u
MM19 a2n a1n a2n VDD pch_mac l=0.03u w=0.17u
MM15 zb a1n net0184 VDD pch_mac l=0.03u w=0.17u
MM14 net0184 a2n VDD VDD pch_mac l=0.03u w=0.17u
MM7 Z zb VDD VDD pch_mac l=0.03u w=0.17u 
MM7_2 Z zb VDD VDD pch_mac l=0.03u w=0.17u 
MM9 a1n A1 VDD VDD pch_mac l=0.03u w=0.17u
.ENDS
.SUBCKT ISOHID2 ISO I Z VDD VSS
MM9 net6 I VSS VSS nch_mac l=30n w=0.14u
MM8 net6 ISO VSS VSS nch_mac l=30n w=0.14u
MM0 Z net6 VSS VSS nch_mac l=30n w=0.14u 
MM0_2 Z net6 VSS VSS nch_mac l=30n w=0.14u 
MM7 net25 ISO VDD VDD pch_mac l=30n w=0.17u
MM3 net6 I net25 VDD pch_mac l=30n w=0.17u
MM1 Z net6 VDD VDD pch_mac l=30n w=0.17u 
MM1_2 Z net6 VDD VDD pch_mac l=30n w=0.17u 
.ENDS
.SUBCKT ISOLOD2 ISO I Z VDD VSS
MM3 net050 ISO VSS VSS nch_mac l=30n w=0.14u
MM9 net14 net050 VSS VSS nch_mac l=30n w=0.14u
MM8 net26 I net14 VSS nch_mac l=30n w=0.14u
MM5 Z net26 VSS VSS nch_mac l=30n w=0.14u 
MM5_2 Z net26 VSS VSS nch_mac l=30n w=0.14u 
MM2 net050 ISO VDD VDD pch_mac l=30n w=0.17u
MM6 net26 I VDD VDD pch_mac l=30n w=170.0n
MM7 net26 net050 VDD VDD pch_mac l=30n w=0.17u
MM4 Z net26 VDD VDD pch_mac l=30n w=0.17u 
MM4_2 Z net26 VDD VDD pch_mac l=30n w=0.17u 
.ENDS
.SUBCKT ISOSRHID2 ISO I Z VDD VDDS VSS
MM7 net36 ISO VDDS VDDS pch_mac l=30.0n w=0.17u
MM1 Z net50 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM1_2 Z net50 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM3 net50 I net36 VDDS pch_mac l=30.0n w=0.17u
MM0 Z net50 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net50 VSS VSS nch_mac l=30.0n w=0.14u 
MM9 net50 I VSS VSS nch_mac l=30.0n w=0.14u
MM8 net50 ISO VSS VSS nch_mac l=30.0n w=0.14u
.ENDS
.SUBCKT ISOSRLOD2 ISO I Z VDD VDDS VSS
MM3 net7 ISO VSS VSS nch_mac l=30.0n w=0.14u
MM9 net11 net7 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net30 I net11 VSS nch_mac l=30.0n w=0.14u
MM5 Z net30 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net30 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 net7 ISO VDDS VDDS pch_mac l=30.0n w=0.17u
MM6 net30 I VDDS VDDS pch_mac l=30.0n w=170n
MM7 net30 net7 VDDS VDDS pch_mac l=30.0n w=0.17u
MM4 Z net30 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM4_2 Z net30 VDDS VDDS pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT LVLHLCD2 I NSLEEP Z VDD VSS
MM1 net0103 I VSS VSS nch_mac l=30.0n w=0.14u
MM4 net084 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u
MM5 Z net0103 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net0103 VSS VSS nch_mac l=30.0n w=0.14u 
MM0 net0103 net084 VSS VSS nch_mac l=30.0n w=0.14u
MM11 net0103 I net069 VDD pch_mac l=30.0n w=0.17u
MM12 net084 NSLEEP VDD VDD pch_mac l=30.0n w=0.17u
MM13 Z net0103 VDD VDD pch_mac l=30.0n w=0.17u 
MM13_2 Z net0103 VDD VDD pch_mac l=30.0n w=0.17u 
MM7 net069 net084 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LVLHLCLOD2 I NSLEEP Z VDD VSS
MM8 Z net28 VSS VSS nch_mac l=30.0n w=0.14u 
MM8_2 Z net28 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 net32 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u
MM3 net28 I net32 VSS nch_mac l=30.0n w=0.14u
MM9 Z net28 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_2 Z net28 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 net28 I VDD VDD pch_mac l=30.0n w=170.0n
MM7 net28 NSLEEP VDD VDD pch_mac l=30.0n w=0.17u
.ENDS
.SUBCKT LVLHLD2 I Z VDD VSS
MM5 net8 I VSS VSS nch_mac l=30.0n w=0.14u
MM0 Z net8 VSS VSS nch_mac l=30.0n w=0.14u 
MM0_2 Z net8 VSS VSS nch_mac l=30.0n w=0.14u 
MM4 net8 I VDD VDD pch_mac l=30.0n w=0.17u
MM1 Z net8 VDD VDD pch_mac l=30.0n w=0.17u 
MM1_2 Z net8 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT LVLLHCD2 I NSLEEP Z VDD VDDL VSS
MM10 N2 N0 N5 VSS nch_mac l=30.0n w=0.14u
MM15 N3 I N5 VSS nch_mac l=30.0n w=0.14u
MM12 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_3 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_4 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM5 Z N3 N5 VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z N3 N5 VSS nch_mac l=30.0n w=0.14u 
MM2 N0 I N5 VSS nch_mac l=30.0n w=0.14u
MM17 N3 I N4 VDD pch_mac l=30.0n w=0.17u 
MM17_2 N3 I N4 VDD pch_mac l=30.0n w=0.17u 
MM17_3 N3 I N4 VDD pch_mac l=30.0n w=0.17u 
MM14 N0 I VDDL VDDL pch_mac l=30.0n w=170.0n
MM16 N2 N0 N1 VDD pch_mac l=30.0n w=0.120u
MM0 Z NSLEEP VDD VDD pch_mac l=30.0n w=0.17u
MM4 Z N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM9 N1 N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_2 N1 N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_3 N1 N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 N4 N2 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 N4 N2 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_3 N4 N2 VDD VDD pch_mac l=30.0n w=0.17u 
.ENDS
.SUBCKT LVLLHCLOD2 I NSLEEP Z VDD VDDL VSS
MM33 N5 N3 N6 VSS nch_mac l=30.0n w=0.14u
MM27 N6 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM27_2 N6 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM27_3 N6 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM27_4 N6 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM28 N3 I N6 VSS nch_mac l=30.0n w=0.14u
MM29 N2 N0 N6 VSS nch_mac l=30.0n w=0.14u
MM30 N0 I N6 VSS nch_mac l=30.0n w=140.0n
MM17 N7 N5 N8 VSS nch_mac l=30.0n w=0.14u
MM32 N8 NSLEEP N6 VSS nch_mac l=30.0n w=0.14u
MM19 Z N7 VSS VSS nch_mac l=30.0n w=0.14u 
MM19_2 Z N7 VSS VSS nch_mac l=30.0n w=0.14u 
MM16 N7 N5 VDD VDD pch_mac l=30.0n w=0.17u
MM15 N7 NSLEEP VDD VDD pch_mac l=30.0n w=0.17u
MM20 Z N7 VDD VDD pch_mac l=30.0n w=0.17u 
MM20_2 Z N7 VDD VDD pch_mac l=30.0n w=0.17u 
MM31 N5 N3 VDD VDD pch_mac l=30.0n w=0.17u
MM21 N0 I VDDL VDDL pch_mac l=30.0n w=0.17u
MM22 N3 I N4 VDD pch_mac l=30.0n w=0.17u 
MM22_2 N3 I N4 VDD pch_mac l=30.0n w=0.17u 
MM22_3 N3 I N4 VDD pch_mac l=30.0n w=0.17u 
MM24 N1 N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM24_2 N1 N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM24_3 N1 N3 VDD VDD pch_mac l=30.0n w=0.17u 
MM25 N4 N2 VDD VDD pch_mac l=30.0n w=0.17u 
MM25_2 N4 N2 VDD VDD pch_mac l=30.0n w=0.17u 
MM25_3 N4 N2 VDD VDD pch_mac l=30.0n w=0.17u 
MM26 N2 N0 N1 VDD pch_mac l=30.0n w=0.120u
.ENDS
.SUBCKT LVLLHD2 I Z VDD VDDL VSS
MM15 net46 I VSS VSS nch_mac l=30.0n w=0.14u
MM10 net64 net57 VSS VSS nch_mac l=30.0n w=0.14u
MM5 Z net46 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net46 VSS VSS nch_mac l=30.0n w=0.14u 
MM2 net57 I VSS VSS nch_mac l=30.0n w=0.14u
MM14 net57 I VDDL VDDL pch_mac l=30.0n w=170.0n
MM4 Z net46 VDD VDD pch_mac l=30.0n w=0.17u 
MM4_2 Z net46 VDD VDD pch_mac l=30.0n w=0.17u 
MM6 net49 net64 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_2 net49 net64 VDD VDD pch_mac l=30.0n w=0.17u 
MM6_3 net49 net64 VDD VDD pch_mac l=30.0n w=0.17u 
MM17 net46 I net49 VDD pch_mac l=30.0n w=0.17u 
MM17_2 net46 I net49 VDD pch_mac l=30.0n w=0.17u 
MM17_3 net46 I net49 VDD pch_mac l=30.0n w=0.17u 
MM9 net44 net46 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_2 net44 net46 VDD VDD pch_mac l=30.0n w=0.17u 
MM9_3 net44 net46 VDD VDD pch_mac l=30.0n w=0.17u 
MM16 net64 net57 net44 VDD pch_mac l=30.0n w=0.120u
.ENDS
.SUBCKT LVLSRLHCD2 I NSLEEP Z VDD VDDS VSS
MM6 N4 N2 VDDS VDDS pch_mac l=30.0n w=170n
MM9 N1 N3 VDDS VDDS pch_mac l=30.0n w=0.12u
MM4 Z N3 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM4_2 Z N3 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM0 Z NSLEEP VDDS VDDS pch_mac l=30.0n w=0.17u
MM16 N2 N0 N1 VDDS pch_mac l=30.0n w=0.12u
MM14 N0 I VDD VDD pch_mac l=30.0n w=170n
MM17 N3 I N4 VDDS pch_mac l=30.0n w=0.17u
MM2 N0 I N5 VSS nch_mac l=30.0n w=0.14u
MM5 Z N3 N5 VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z N3 N5 VSS nch_mac l=30.0n w=0.14u 
MM12 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_2 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_3 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_4 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM12_5 N5 NSLEEP VSS VSS nch_mac l=30.0n w=0.14u 
MM15 N3 I N5 VSS nch_mac l=30.0n w=0.14u 
MM15_2 N3 I N5 VSS nch_mac l=30.0n w=0.14u 
MM15_3 N3 I N5 VSS nch_mac l=30.0n w=0.14u 
MM10 N2 N0 N5 VSS nch_mac l=30.0n w=0.14u 
MM10_2 N2 N0 N5 VSS nch_mac l=30.0n w=0.14u 
MM10_3 N2 N0 N5 VSS nch_mac l=30.0n w=0.14u 
.ENDS
.SUBCKT LVLSRLHD2 I Z VDD VDDS VSS
MM16 net39 net31 net9 VDDS pch_mac l=30.0n w=0.12u
MM9 net9 net11 VDDS VDDS pch_mac l=30.0n w=0.12u
MM17 net11 I net17 VDDS pch_mac l=30.0n w=0.17u
MM6 net17 net39 VDDS VDDS pch_mac l=30.0n w=170n
MM4 Z net11 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM4_2 Z net11 VDDS VDDS pch_mac l=30.0n w=0.17u 
MM14 net31 I VDD VDD pch_mac l=30.0n w=170n
MM2 net31 I VSS VSS nch_mac l=30.0n w=0.14u
MM5 Z net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM5_2 Z net11 VSS VSS nch_mac l=30.0n w=0.14u 
MM10 net39 net31 VSS VSS nch_mac l=30.0n w=0.14u 
MM10_2 net39 net31 VSS VSS nch_mac l=30.0n w=0.14u 
MM10_3 net39 net31 VSS VSS nch_mac l=30.0n w=0.14u 
MM15 net11 I VSS VSS nch_mac l=30.0n w=0.14u 
MM15_2 net11 I VSS VSS nch_mac l=30.0n w=0.14u 
MM15_3 net11 I VSS VSS nch_mac l=30.0n w=0.14u 
.ENDS
.SUBCKT AD1V4 A B CI CO S VDD VSS
MM24 S net181 VDD VDD pch_mac W=400.00n L=30.00n
MM16 net181 CI net152 VDD pch_mac W=200.00n L=30.00n
MM14 net144 B VDD VDD pch_mac W=200.00n L=30.00n
MM15 net152 A net144 VDD pch_mac W=200.00n L=30.00n
MM13 net181 net177 net129 VDD pch_mac W=200.00n L=30.00n
MM12 net129 CI VDD VDD pch_mac W=200.00n L=30.00n
MM10 net129 B VDD VDD pch_mac W=200.00n L=30.00n
MM11 net129 A VDD VDD pch_mac W=200.00n L=30.00n
MM7 net177 A net124 VDD pch_mac W=200.00n L=30.00n
MM6 net124 B VDD VDD pch_mac W=200.00n L=30.00n
MM5 CO net177 VDD VDD pch_mac W=400.00n L=30.00n
MM1 net177 CI net101 VDD pch_mac W=200.00n L=30.00n
MM0 net101 B VDD VDD pch_mac W=200.00n L=30.00n
MM28 net101 A VDD VDD pch_mac W=200.00n L=30.00n
MM25 S net181 VSS VSS nch_mac W=400.00n L=30.00n
MM23 net189 CI VSS VSS nch_mac W=175.00n L=30.00n
MM20 net197 B VSS VSS nch_mac W=200.00n L=30.00n
MM19 net193 A net197 VSS nch_mac W=200.00n L=30.00n
MM21 net189 A VSS VSS nch_mac W=200.00n L=30.00n
MM18 net181 CI net193 VSS nch_mac W=175.00n L=30.00n
MM17 net181 net177 net189 VSS nch_mac W=175.00n L=30.00n
MM9 net177 A net173 VSS nch_mac W=200.00n L=30.00n
MM8 net173 B VSS VSS nch_mac W=200.00n L=30.00n
MM4 CO net177 VSS VSS nch_mac W=400.00n L=30.00n
MM3 net177 CI net157 VSS nch_mac W=200.00n L=30.00n
MM2 net157 B VSS VSS nch_mac W=200.00n L=30.00n
MM29 net157 A VSS VSS nch_mac W=200.00n L=30.00n
MM22 net189 B VSS VSS nch_mac W=200.00n L=30.00n
.ENDS AD1V4
.SUBCKT ADH1V4 A B CO S VDD VSS
MM5 CO nandab VDD VDD pch_mac W=400.00n L=30.00n
MM3 S net121 VDD VDD pch_mac W=400.00n L=30.00n
MM1 net121 nandab VDD VDD pch_mac W=200.00n L=30.00n
MM7 net121 A net96 VDD pch_mac W=200.00n L=30.00n
MM0 nandab B VDD VDD pch_mac W=200.00n L=30.00n
MM28 nandab A VDD VDD pch_mac W=200.00n L=30.00n
MM6 net96 B VDD VDD pch_mac W=200.00n L=30.00n
MM2 net129 B VSS VSS nch_mac W=200.00n L=30.00n
MM29 net129 A VSS VSS nch_mac W=200.00n L=30.00n
MM8 net125 B VSS VSS nch_mac W=200.00n L=30.00n
MM10 net121 nandab net129 VSS nch_mac W=200.00n L=30.00n
MM9 nandab A net125 VSS nch_mac W=200.00n L=30.00n
MM11 S net121 VSS VSS nch_mac W=400.00n L=30.00n
MM4 CO nandab VSS VSS nch_mac W=400.00n L=30.00n
.ENDS ADH1V4
.SUBCKT AND2V4 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VSS nch_mac W=0.2u L=30.00n
MM2 Z net11 VSS VSS nch_mac W=0.4u L=30.00n
MMN1 net18 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM3 Z net11 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net11 A2 VDD VDD pch_mac W=0.2u L=30.00n
MMP1 net11 A1 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS AND2V4
.SUBCKT AND3V4 A1 A2 A3 Z VDD VSS
MM1 net11 A1 net18 VSS nch_mac W=0.2u L=30.00n
MM2 Z net11 VSS VSS nch_mac W=0.4u L=30.00n
MM4 net_043 A3 VSS VSS nch_mac W=0.2u L=30.00n
MMN1 net18 A2 net_043 VSS nch_mac W=0.2u L=30.00n
MM5 net11 A3 VDD VDD pch_mac W=0.2u L=30.00n
MM3 Z net11 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net11 A2 VDD VDD pch_mac W=0.2u L=30.00n
MMP1 net11 A1 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS AND3V4
.SUBCKT AND4V4 A1 A2 A3 A4 Z VDD VSS
MM6 net_042 A4 VSS VSS nch_mac W=0.2u L=30.00n
MM1 net11 A1 net18 VSS nch_mac W=0.2u L=30.00n
MM2 Z net11 VSS VSS nch_mac W=0.4u L=30.00n
MM4 net_054 A3 net_042 VSS nch_mac W=0.2u L=30.00n
MMN1 net18 A2 net_054 VSS nch_mac W=0.2u L=30.00n
MM7 net11 A4 VDD VDD pch_mac W=0.2u L=30.00n
MM5 net11 A3 VDD VDD pch_mac W=0.2u L=30.00n
MM3 Z net11 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net11 A2 VDD VDD pch_mac W=0.2u L=30.00n
MMP1 net11 A1 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS AND4V4
.SUBCKT AO112V4 A1 A2 B C Z VDD VSS
MM5 Z net6 VSS VSS nch_mac W=0.4u L=30.00n
MM8 net30 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM9 net6 A1 net30 VSS nch_mac W=0.2u L=30.00n
MM3 net6 B VSS VSS nch_mac W=0.2u L=30.00n
MM4 net6 C VSS VSS nch_mac W=0.2u L=30.00n
MM28 net6 A1 net056 VDD pch_mac W=0.2u L=30.00n
MM0 net6 A2 net056 VDD pch_mac W=0.2u L=30.00n
MM1 net21 C VDD VDD pch_mac W=0.2u L=30.00n
MM2 net056 B net21 VDD pch_mac W=0.2u L=30.00n
MM6 Z net6 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS AO112V4
.SUBCKT AO12V4 A1 A2 B Z VDD VSS
MM4 Z net048 VSS VSS nch_mac W=0.4u L=30.00n
MM2 net048 B VSS VSS nch_mac W=0.2u L=30.00n
MM9 net048 A1 net13 VSS nch_mac W=0.2u L=30.00n
MM8 net13 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM3 Z net048 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net043 B VDD VDD pch_mac W=0.2u L=30.00n
MM0 net048 A2 net043 VDD pch_mac W=0.2u L=30.00n
MM28 net048 A1 net043 VDD pch_mac W=0.2u L=30.00n
.ENDS AO12V4
.SUBCKT AO13V4 A1 A2 A3 B Z VDD VSS
MM5 Z net34 VDD VDD pch_mac W=0.4u L=30.00n
MM4 net34 A3 net37 VDD pch_mac W=0.2u L=30.00n
MM0 net34 A2 net37 VDD pch_mac W=0.2u L=30.00n
MM28 net34 A1 net37 VDD pch_mac W=0.2u L=30.00n
MM1 net37 B VDD VDD pch_mac W=0.2u L=30.00n
MM8 net50 A2 net42 VSS nch_mac W=0.2u L=30.00n
MM6 Z net34 VSS VSS nch_mac W=0.4u L=30.00n
MM9 net34 A1 net50 VSS nch_mac W=0.2u L=30.00n
MM3 net42 A3 VSS VSS nch_mac W=0.2u L=30.00n
MM2 net34 B VSS VSS nch_mac W=0.2u L=30.00n
.ENDS AO13V4
.SUBCKT AO1B2V4 A1 A2 B Z VDD VSS
MM2 Z B net030 VSS nch_mac W=0.4u L=30.00n
MM3 net030 net055 VSS VSS nch_mac W=0.4u L=30.00n
MM1 net055 A1 net18 VSS nch_mac W=0.175u L=30.00n
MMN1 net18 A2 VSS VSS nch_mac W=0.175u L=30.00n
MM4 Z net055 VDD VDD pch_mac W=0.4u L=30.00n
MM5 Z B VDD VDD pch_mac W=0.35u L=30.00n
MM0 net055 A2 VDD VDD pch_mac W=0.175u L=30.00n
MMP1 net055 A1 VDD VDD pch_mac W=0.175u L=30.00n
.ENDS AO1B2V4
.SUBCKT AO212V4 A1 A2 B1 B2 C Z VDD VSS
MM0 net36 B2 VDD VDD pch_mac W=0.2u L=30.00n
MM28 net36 B1 VDD VDD pch_mac W=0.2u L=30.00n
MM6 net48 A1 net43 VDD pch_mac W=0.2u L=30.00n
MM1 net43 C net36 VDD pch_mac W=0.2u L=30.00n
MM10 Z net48 VDD VDD pch_mac W=0.4u L=30.00n
MM5 net48 A2 net43 VDD pch_mac W=0.2u L=30.00n
MM7 Z net48 VSS VSS nch_mac W=400.00n L=30.00n
MM8 net60 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM3 net68 B2 VSS VSS nch_mac W=0.2u L=30.00n
MM9 net48 A1 net60 VSS nch_mac W=0.2u L=30.00n
MM2 net48 B1 net68 VSS nch_mac W=0.2u L=30.00n
MM4 net48 C VSS VSS nch_mac W=0.2u L=30.00n
.ENDS AO212V4
.SUBCKT AO222V4 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM12 Z net81 VDD VDD pch_mac W=0.4u L=30.00n
MM10 net81 A2 net48 VDD pch_mac W=0.175u L=30.00n
MM28 net48 B1 net40 VDD pch_mac W=0.175u L=30.00n
MM0 net48 B2 net40 VDD pch_mac W=0.175u L=30.00n
MM1 net81 A1 net48 VDD pch_mac W=0.175u L=30.00n
MM6 net40 C1 VDD VDD pch_mac W=0.175u L=30.00n
MM5 net40 C2 VDD VDD pch_mac W=0.175u L=30.00n
MM11 Z net81 VSS VSS nch_mac W=0.4u L=30.00n
MM7 net61 C2 VSS VSS nch_mac W=0.19u L=30.00n
MM3 net65 B2 VSS VSS nch_mac W=0.19u L=30.00n
MM4 net81 C1 net61 VSS nch_mac W=0.19u L=30.00n
MM2 net81 B1 net65 VSS nch_mac W=0.19u L=30.00n
MM9 net81 A1 net69 VSS nch_mac W=0.19u L=30.00n
MM8 net69 A2 VSS VSS nch_mac W=0.19u L=30.00n
.ENDS AO222V4
.SUBCKT AO22V4 A1 A2 B1 B2 Z VDD VSS
MM1 net48 A1 net35 VDD pch_mac W=0.2u L=30.00n
MM5 Z net48 VDD VDD pch_mac W=0.4u L=30.00n
MM2 net48 A2 net35 VDD pch_mac W=0.2u L=30.00n
MM0 net35 B2 VDD VDD pch_mac W=0.2u L=30.00n
MM28 net35 B1 VDD VDD pch_mac W=0.2u L=30.00n
MM8 net44 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM6 Z net48 VSS VSS nch_mac W=0.4u L=30.00n
MM3 net48 B1 net56 VSS nch_mac W=0.2u L=30.00n
MM9 net48 A1 net44 VSS nch_mac W=0.2u L=30.00n
MM4 net56 B2 VSS VSS nch_mac W=0.2u L=30.00n
.ENDS AO22V4
.SUBCKT AO32V4 A1 A2 A3 B1 B2 Z VDD VSS
MM3 net31 A3 VSS VSS nch_mac W=200.0n L=30.00n
MM2 net35 B1 net47 VSS nch_mac W=200.0n L=30.00n
MM9 net35 A1 net43 VSS nch_mac W=200.0n L=30.00n
MM8 net43 A2 net31 VSS nch_mac W=200.0n L=30.00n
MM5 net47 B2 VSS VSS nch_mac W=200.0n L=30.00n
MM7 Z net35 VSS VSS nch_mac W=400.0n L=30.00n
MM28 net7 A1 VDD VDD pch_mac W=200.0n L=30.00n
MM4 net7 A3 VDD VDD pch_mac W=200.0n L=30.00n
MM0 net7 A2 VDD VDD pch_mac W=200.0n L=30.00n
MM1 net35 B2 net7 VDD pch_mac W=200.0n L=30.00n
MM6 net35 B1 net7 VDD pch_mac W=200.0n L=30.00n
MM10 Z net35 VDD VDD pch_mac W=400.0n L=30.00n
.ENDS AO32V4
.SUBCKT AO33V4 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM2 net40 B1 net20 VSS nch_mac W=0.2u L=30.00n
MM9 net40 A1 net16 VSS nch_mac W=0.2u L=30.00n
MM8 net16 A2 net28 VSS nch_mac W=0.2u L=30.00n
MM5 net20 B2 net24 VSS nch_mac W=0.2u L=30.00n
MM11 net24 B3 VSS VSS nch_mac W=0.2u L=30.00n
MM3 net28 A3 VSS VSS nch_mac W=0.2u L=30.00n
MM7 Z net40 VSS VSS nch_mac W=0.4u L=30.00n
MM1 net40 A2 net43 VDD pch_mac W=0.2u L=30.00n
MM6 net40 A1 net43 VDD pch_mac W=0.2u L=30.00n
MM12 net40 A3 net43 VDD pch_mac W=0.2u L=30.00n
MM10 Z net40 VDD VDD pch_mac W=0.4u L=30.00n
MM28 net43 B1 VDD VDD pch_mac W=0.2u L=30.00n
MM4 net43 B3 VDD VDD pch_mac W=0.2u L=30.00n
MM0 net43 B2 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS AO33V4
.SUBCKT AOI112V4 A1 A2 B C ZN VDD VSS
MMP1 net_58 B net2 VDD pch_mac W=0.4u L=30.00n
MM0 net2 C VDD VDD pch_mac W=0.4u L=30.00n
MM5 ZN A2 net_58 VDD pch_mac W=0.4u L=30.00n
MM7 ZN A1 net_58 VDD pch_mac W=0.4u L=30.00n
MM1 ZN A1 net4 VSS nch_mac W=0.4u L=30.00n
MMN1 net4 A2 VSS VSS nch_mac W=0.4u L=30.00n
MM4 ZN B VSS VSS nch_mac W=0.4u L=30.00n
MM6 ZN C VSS VSS nch_mac W=0.4u L=30.00n
.ENDS AOI112V4
.SUBCKT AOI12V4 A1 A2 B ZN VDD VSS
MM7 ZN A1 net_37 VDD pch_mac W=0.4u L=30.00n
MM5 ZN A2 net_37 VDD pch_mac W=0.4u L=30.00n
MM0 net_37 B VDD VDD pch_mac W=0.4u L=30.00n
MMN1 net4 A2 VSS VSS nch_mac W=0.4u L=30.00n
MM6 ZN B VSS VSS nch_mac W=0.4u L=30.00n
MM1 ZN A1 net4 VSS nch_mac W=0.4u L=30.00n
.ENDS AOI12V4
.SUBCKT AOI13V4 A1 A2 A3 B ZN VDD VSS
MM9 ZN A1 net45 VSS nch_mac W=0.4u L=30.00n
MM8 net45 A2 net53 VSS nch_mac W=0.4u L=30.00n
MM2 ZN B VSS VSS nch_mac W=0.4u L=30.00n
MM3 net53 A3 VSS VSS nch_mac W=0.4u L=30.00n
MM0 ZN A2 net64 VDD pch_mac W=0.4u L=30.00n
MM28 ZN A1 net64 VDD pch_mac W=0.4u L=30.00n
MM4 ZN A3 net64 VDD pch_mac W=0.4u L=30.00n
MM1 net64 B VDD VDD pch_mac W=0.4u L=30.00n
.ENDS AOI13V4
.SUBCKT AOI212V4 A1 A2 B1 B2 C ZN VDD VSS
MM7 net53 B1 VDD VDD pch_mac W=0.4u L=30.00n
MM8 ZN A2 net72 VDD pch_mac W=0.4u L=30.00n
MM5 net53 B2 VDD VDD pch_mac W=0.4u L=30.00n
MM0 ZN A1 net72 VDD pch_mac W=0.4u L=30.00n
MMP1 net72 C net53 VDD pch_mac W=0.4u L=30.00n
MMN1 net81 A2 VSS VSS nch_mac W=0.4u L=30.00n
MM6 ZN C VSS VSS nch_mac W=0.4u L=30.00n
MM4 ZN B1 N3 VSS nch_mac W=0.4u L=30.00n
MM9 N3 B2 VSS VSS nch_mac W=0.4u L=30.00n
MM1 ZN A1 net81 VSS nch_mac W=0.4u L=30.00n
.ENDS AOI212V4
.SUBCKT AOI21BV4 A B1 B2 ZN VDD VSS
MM3 net21 A VSS VSS nch_mac W=0.175u L=30.00n
MM2 ZN net21 VSS VSS nch_mac W=0.4u L=30.00n
MM9 ZN B1 net33 VSS nch_mac W=0.4u L=30.00n
MM8 net33 B2 VSS VSS nch_mac W=0.4u L=30.00n
MM4 net21 A VDD VDD pch_mac W=0.175u L=30.00n
MM1 ZN net21 net17 VDD pch_mac W=0.4u L=30.00n
MM0 net17 B2 VDD VDD pch_mac W=0.4u L=30.00n
MM28 net17 B1 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS AOI21BV4
.SUBCKT AOI222V4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM6 ZN C1 net4 VSS nch_mac W=0.4u L=30.00n
MM10 net4 C2 VSS VSS nch_mac W=0.4u L=30.00n
MM9 net5 B2 VSS VSS nch_mac W=0.4u L=30.00n
MM1 ZN A1 net6 VSS nch_mac W=0.4u L=30.00n
MM4 ZN B1 net5 VSS nch_mac W=0.4u L=30.00n
MMN1 net6 A2 VSS VSS nch_mac W=0.4u L=30.00n
MM8 net2 B2 net1 VDD pch_mac W=0.4u L=30.00n
MM11 ZN A2 net2 VDD pch_mac W=0.4u L=30.00n
MM7 net1 C1 VDD VDD pch_mac W=0.4u L=30.00n
MM5 net1 C2 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net2 B1 net1 VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 net2 VDD pch_mac W=0.4u L=30.00n
.ENDS AOI222V4
.SUBCKT AOI22BBV4 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 A1 VSS VSS nch_mac W=0.175u L=30.00n
MM2 net24 A2 VSS VSS nch_mac W=0.175u L=30.00n
MM0 ZN B1 net050 VSS nch_mac W=0.435u L=30.00n
MM7 net050 B2 VSS VSS nch_mac W=0.4u L=30.00n
MMN1 ZN net24 VSS VSS nch_mac W=0.4u L=30.00n
MM6 ZN B2 net078 VDD pch_mac W=0.4u L=30.00n
MM4 net24 A1 net074 VDD pch_mac W=0.175u L=30.00n
MM5 net074 A2 VDD VDD pch_mac W=0.175u L=30.00n
MM1 net078 net24 VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN B1 net078 VDD pch_mac W=0.435u L=30.00n
.ENDS AOI22BBV4
.SUBCKT AOI22V4 A1 A2 B1 B2 ZN VDD VSS
MM5 N69 B2 VDD VDD pch_mac W=0.4u L=30.00n
MM7 N69 B1 VDD VDD pch_mac W=0.4u L=30.00n
MM0 ZN A1 N69 VDD pch_mac W=0.4u L=30.00n
MM8 ZN A2 N69 VDD pch_mac W=0.4u L=30.00n
MM1 ZN A1 N49 VSS nch_mac W=0.4u L=30.00n
MM9 N64 B2 VSS VSS nch_mac W=0.4u L=30.00n
MM4 ZN B1 N64 VSS nch_mac W=0.4u L=30.00n
MMN1 N49 A2 VSS VSS nch_mac W=0.4u L=30.00n
.ENDS AOI22V4
.SUBCKT AOI32V4 A1 A2 A3 B1 B2 ZN VDD VSS
MM6 ZN B1 net5 VSS nch_mac W=400.00n L=30.00n
MM1 ZN A1 net3 VSS nch_mac W=400.00n L=30.00n
MM9 net4 A3 VSS VSS nch_mac W=400.00n L=30.00n
MM11 net5 B2 VSS VSS nch_mac W=400.00n L=30.00n
MMN1 net3 A2 net4 VSS nch_mac W=400.00n L=30.00n
MM8 net1 A3 VDD VDD pch_mac W=400.00n L=30.00n
MM10 ZN B2 net1 VDD pch_mac W=400.00n L=30.00n
MM7 net1 A1 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net1 A2 VDD VDD pch_mac W=400.00n L=30.00n
MM0 ZN B1 net1 VDD pch_mac W=400.00n L=30.00n
.ENDS AOI32V4
.SUBCKT AOI33V4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM12 net_69 B3 VSS VSS nch_mac W=400.00n L=30.00n
MM6 ZN B1 net5 VSS nch_mac W=400.00n L=30.00n
MM1 ZN A1 net3 VSS nch_mac W=400.00n L=30.00n
MM9 net4 A3 VSS VSS nch_mac W=400.00n L=30.00n
MM11 net5 B2 net_69 VSS nch_mac W=400.00n L=30.00n
MMN1 net3 A2 net4 VSS nch_mac W=400.00n L=30.00n
MM8 net1 A3 VDD VDD pch_mac W=400.00n L=30.00n
MM10 ZN B2 net1 VDD pch_mac W=400.00n L=30.00n
MM7 net1 A1 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net1 A2 VDD VDD pch_mac W=400.00n L=30.00n
MM13 ZN B3 net1 VDD pch_mac W=400.00n L=30.00n
MM0 ZN B1 net1 VDD pch_mac W=400.00n L=30.00n
.ENDS AOI33V4
.SUBCKT BUFV4 I Z VDD VSS
MM1 Z net25 VSS VSS nch_mac W=0.4u L=30.00n
MM2 net25 I VSS VSS nch_mac W=0.2u L=30.00n
MM0 Z net25 VDD VDD pch_mac W=0.4u L=30.00n
MM3 net25 I VDD VDD pch_mac W=0.2u L=30.00n
.ENDS BUFV4
.SUBCKT CLKAND2V4 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VSS nch_mac W=0.2u L=30.00n
MM2 Z net11 VSS VSS nch_mac W=0.24u L=30.00n
MMN1 net18 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM3 Z net11 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net11 A2 VDD VDD pch_mac W=0.2u L=30.00n
MMP1 net11 A1 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS CLKAND2V4
.SUBCKT CLKBUFV4 I Z VDD VSS
MM1 Z net25 VSS VSS nch_mac W=0.24u L=30.00n
MM2 net25 I VSS VSS nch_mac W=0.12u L=30.00n
MM0 Z net25 VDD VDD pch_mac W=0.4u L=30.00n
MM3 net25 I VDD VDD pch_mac W=0.2u L=30.00n
.ENDS CLKBUFV4
.SUBCKT CLKINV4 I ZN VDD VSS
MM2 ZN I VSS VSS nch_mac W=0.24u L=30.00n
MM3 ZN I VDD VDD pch_mac W=0.4u L=30.00n
.ENDS CLKINV4
.SUBCKT CLKLAHAQV4 CK E Q TE VDD VSS
MM12 s ten net217 VDD pch_mac W=0.2u L=30.00n
MM14 net217 c VDD VDD pch_mac W=0.2u L=30.00n
MM13 s pm net217 VDD pch_mac W=0.2u L=30.00n
MM15 Q s VDD VDD pch_mac W=0.4u L=30.00n
MM22 nt13 m VDD VDD pch_mac W=0.125u L=30.00n
MM23 pm c nt13 VDD pch_mac W=0.125u L=30.00n
MM16 nt11 cn VDD VDD pch_mac W=0.125u L=30.00n
MM17 pm E nt11 VDD pch_mac W=0.125u L=30.00n
MM21 m pm VDD VDD pch_mac W=0.125u L=30.00n
MM19 c cn VDD VDD pch_mac W=0.125u L=30.00n
MM20 ten TE VDD VDD pch_mac W=0.125u L=30.00n
MM18 cn CK VDD VDD pch_mac W=0.125u L=30.00n
MM7 Q s VSS VSS nch_mac W=0.24u L=30.00n
MM9 nt22 ten VSS VSS nch_mac W=120.00n L=30.00n
MM1 nt12 E VSS VSS nch_mac W=0.125u L=30.00n
MM8 s c VSS VSS nch_mac W=120.00n L=30.00n
MM0 pm c nt12 VSS nch_mac W=0.125u L=30.00n
MM6 s pm nt22 VSS nch_mac W=120.00n L=30.00n
MM11 nt14 cn VSS VSS nch_mac W=0.125u L=30.00n
MM5 ten TE VSS VSS nch_mac W=0.125u L=30.00n
MM10 pm m nt14 VSS nch_mac W=0.125u L=30.00n
MM3 cn CK VSS VSS nch_mac W=0.125u L=30.00n
MM4 c cn VSS VSS nch_mac W=0.125u L=30.00n
MM2 m pm VSS VSS nch_mac W=0.125u L=30.00n
.ENDS CLKLAHAQV4
.SUBCKT CLKLAHQV4 CK E Q TE VDD VSS
MM9 hnet21 m VDD VDD pch_mac W=120.00n L=30.00n
MM5 m pm VDD VDD pch_mac W=120.00n L=30.00n
MM2 hnet13 cn VDD VDD pch_mac W=0.125u L=30.00n
MM4 pm E hnet11 VDD pch_mac W=0.15u L=30.00n
MM10 pm c hnet21 VDD pch_mac W=120.00n L=30.00n
MM3 hnet11 TE hnet13 VDD pch_mac W=0.15u L=30.00n
MM8 Q s VDD VDD pch_mac W=0.4u L=30.00n
MM6 hnet31 pm VDD VDD pch_mac W=0.2u L=30.00n
MM0 cn CK VDD VDD pch_mac W=0.125u L=30.00n
MM7 s c hnet31 VDD pch_mac W=0.2u L=30.00n
MM12 c cn VDD VDD pch_mac W=0.15u L=30.00n
MM21 hnet22 cn VSS VSS nch_mac W=0.125u L=30.00n
MM14 hnet12 E VSS VSS nch_mac W=0.125u L=30.00n
MM20 pm m hnet22 VSS nch_mac W=0.125u L=30.00n
MM13 pm c hnet12 VSS nch_mac W=0.125u L=30.00n
MM15 hnet12 TE VSS VSS nch_mac W=0.125u L=30.00n
MM1 c cn VSS VSS nch_mac W=0.125u L=30.00n
MM11 cn CK VSS VSS nch_mac W=0.125u L=30.00n
MM19 Q s VSS VSS nch_mac W=0.24u L=30.00n
MM16 m pm VSS VSS nch_mac W=120.00n L=30.00n
MM18 s c VSS VSS nch_mac W=120.00n L=30.00n
MM17 s pm VSS VSS nch_mac W=120.00n L=30.00n
.ENDS CLKLAHQV4
.SUBCKT CLKLANAQV4 CK E Q TE VDD VSS
MM15 m pm VDD VDD pch_mac W=0.12u L=30.00n
MM13 nt11 E VDD VDD pch_mac W=0.125u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.125u L=30.00n
MM20 nt13 cn VDD VDD pch_mac W=0.125u L=30.00n
MM14 pm c nt11 VDD pch_mac W=0.125u L=30.00n
MM21 pm m nt13 VDD pch_mac W=0.125u L=30.00n
MM17 s c VDD VDD pch_mac W=0.12u L=30.00n
MM18 s m nt21 VDD pch_mac W=0.12u L=30.00n
MM16 nt21 TE VDD VDD pch_mac W=0.12u L=30.00n
MM19 Q s VDD VDD pch_mac W=0.4u L=30.00n
MM12 c cn VDD VDD pch_mac W=0.125u L=30.00n
MM2 pm E nt12 VSS nch_mac W=0.125u L=30.00n
MM0 cn CK VSS VSS nch_mac W=0.125u L=30.00n
MM4 m pm VSS VSS nch_mac W=0.12u L=30.00n
MM9 pm c nt14 VSS nch_mac W=0.125u L=30.00n
MM10 nt14 m VSS VSS nch_mac W=0.125u L=30.00n
MM1 c cn VSS VSS nch_mac W=0.125u L=30.00n
MM3 nt12 cn VSS VSS nch_mac W=0.125u L=30.00n
MM7 s TE net256 VSS nch_mac W=0.2u L=30.00n
MM8 Q s VSS VSS nch_mac W=0.24u L=30.00n
MM6 s m net256 VSS nch_mac W=0.2u L=30.00n
MM5 net256 c VSS VSS nch_mac W=0.2u L=30.00n
.ENDS CLKLANAQV4
.SUBCKT CLKLANQV4 CK E Q TE VDD VSS
MM10 net220 net196 net151 VDD pch_mac W=120.00n L=30.00n
MM6 net196 net220 VDD VDD pch_mac W=0.12u L=30.00n
MM8 net220 c net163 VDD pch_mac W=0.15u L=30.00n
MM13 net151 cn VDD VDD pch_mac W=120.00n L=30.00n
MM20 net159 TE VDD VDD pch_mac W=0.15u L=30.00n
MM1 net163 E net159 VDD pch_mac W=0.15u L=30.00n
MM18 Q net200 VDD VDD pch_mac W=0.4u L=30.00n
MM5 c cn VDD VDD pch_mac W=0.125u L=30.00n
MM3 cn CK VDD VDD pch_mac W=0.125u L=30.00n
MM14 net200 c VDD VDD pch_mac W=0.2u L=30.00n
MM15 net200 net196 VDD VDD pch_mac W=0.2u L=30.00n
MM19 Q net200 VSS VSS nch_mac W=0.24u L=30.00n
MM9 net228 cn VSS VSS nch_mac W=0.125u L=30.00n
MM4 c cn VSS VSS nch_mac W=0.125u L=30.00n
MM12 net220 c net192 VSS nch_mac W=0.125u L=30.00n
MM17 net200 c net208 VSS nch_mac W=0.165u L=30.00n
MM7 net196 net220 VSS VSS nch_mac W=0.125u L=30.00n
MM0 cn CK VSS VSS nch_mac W=0.125u L=30.00n
MM16 net208 net196 VSS VSS nch_mac W=0.165u L=30.00n
MM21 net220 TE net228 VSS nch_mac W=0.145u L=30.00n
MM2 net220 E net228 VSS nch_mac W=0.145u L=30.00n
MM11 net192 net196 VSS VSS nch_mac W=0.125u L=30.00n
.ENDS CLKLANQV4
.SUBCKT CLKMUX2V4 I0 I1 S Z VDD VSS
MM3 net_52 I0 net077 VSS nch_mac W=200.00n L=30.00n
MM2 net077 SN VSS VSS nch_mac W=200.00n L=30.00n
MM53 SN S VSS VSS nch_mac W=200.0n L=30.00n
MM1 net065 S VSS VSS nch_mac W=200.00n L=30.00n
MM49 net_52 I1 net065 VSS nch_mac W=200.00n L=30.00n
MM51 Z net_52 VSS VSS nch_mac W=240.00n L=30.00n
MM4 net096 S VDD VDD pch_mac W=200.0n L=30.00n
MM5 net_52 SN net096 VDD pch_mac W=200.0n L=30.00n
MM0 net096 I1 VDD VDD pch_mac W=200.0n L=30.00n
MM54 SN S VDD VDD pch_mac W=200.00n L=30.00n
MM52 Z net_52 VDD VDD pch_mac W=400.0n L=30.00n
MM50 net_52 I0 net096 VDD pch_mac W=200.0n L=30.00n
.ENDS CLKMUX2V4
.SUBCKT CLKNAND2V4 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VSS nch_mac W=0.4u L=30.00n
MMN1 net18 A2 VSS VSS nch_mac W=0.4u L=30.00n
MM0 ZN A2 VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS CLKNAND2V4
.SUBCKT CLKNOR2V4 A1 A2 ZN VDD VSS
MMN1 ZN A1 VSS VSS nch_mac W=0.24u L=30.00n
MM0 ZN A2 VSS VSS nch_mac W=0.24u L=30.00n
MMP1 net15 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM1 ZN A1 net15 VDD pch_mac W=0.4u L=30.00n
.ENDS CLKNOR2V4
.SUBCKT CLKOR2V4 A1 A2 Z VDD VSS
MMN1 net12 A1 VSS VSS nch_mac W=120.00n L=30.00n
MM2 Z net12 VSS VSS nch_mac W=0.24u L=30.00n
MM0 net12 A2 VSS VSS nch_mac W=120.00n L=30.00n
MMP1 net23 A2 VDD VDD pch_mac W=0.2u L=30.00n
MM4 Z net12 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net12 A1 net23 VDD pch_mac W=0.2u L=30.00n
.ENDS CLKOR2V4
.SUBCKT CLKXOR2V4 A1 A2 Z VDD VSS
MM0 net73 A2 VSS VSS nch_mac W=200.0n L=30.00n
MMN1 net73 A1 VSS VSS nch_mac W=200.0n L=30.00n
MM9 Z A1 net057 VSS nch_mac W=400.0n L=30.00n
MM4 Z net73 VSS VSS nch_mac W=400.0n L=30.00n
MM3 net057 A2 VSS VSS nch_mac W=400.0n L=30.00n
MM1 net73 A1 net52 VDD pch_mac W=200.0n L=30.00n
MMP1 net52 A2 VDD VDD pch_mac W=200.0n L=30.00n
MM10 Z A1 net048 VDD pch_mac W=400.0n L=30.00n
MM11 Z A2 net048 VDD pch_mac W=400.0n L=30.00n
MM7 net048 net73 VDD VDD pch_mac W=400.0n L=30.00n
.ENDS CLKXOR2V4
.SUBCKT DEL1V4 I Z VDD VSS
MM6 net19 net022 VSS VSS nch_mac W=120.00n L=30.00n
MM1 net022 net11 VSS VSS nch_mac W=120.00n L=30.00n
MM0 Z net19 VSS VSS nch_mac W=400.0n L=30.00n
MM5 net11 I VSS VSS nch_mac W=120.00n L=30.00n
MM7 net19 net022 VDD VDD pch_mac W=200.00n L=30.00n
MM2 net022 net11 VDD VDD pch_mac W=200.00n L=30.00n
MM3 Z net19 VDD VDD pch_mac W=400.00n L=30.00n
MM4 net11 I VDD VDD pch_mac W=200.00n L=30.00n
.ENDS DEL1V4
.SUBCKT DEL2V4 I Z VDD VSS
MM10 net018 I VSS VSS nch_mac W=0.12u L=30.00n
MM6 net026 net018 net022 VSS nch_mac W=120.00n L=30.00n
MM7 net022 net018 VSS VSS nch_mac W=120.00n L=30.00n
MM2 net19 net026 net11 VSS nch_mac W=120.00n L=30.00n
MM0 Z net19 VSS VSS nch_mac W=400.00n L=30.00n
MM5 net11 net026 VSS VSS nch_mac W=120.00n L=30.00n
MM8 net026 net018 net053 VDD pch_mac W=200.0n L=30.00n
MM9 net053 net018 VDD VDD pch_mac W=200.0n L=30.00n
MM11 net018 I VDD VDD pch_mac W=200.0n L=30.00n
MM1 net19 net026 net46 VDD pch_mac W=200.0n L=30.00n
MM3 Z net19 VDD VDD pch_mac W=400.0n L=30.00n
MM4 net46 net026 VDD VDD pch_mac W=200.0n L=30.00n
.ENDS DEL2V4
.SUBCKT DEL4V4 I Z VDD VSS
MM16 net048 net11 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net044 net11 net048 VSS nch_mac W=120.00n L=30.00n
MM18 net040 net23 net036 VSS nch_mac W=120.00n L=30.00n
MM19 net036 net23 VSS VSS nch_mac W=120.00n L=30.00n
MM13 net19 net23 net3 VSS nch_mac W=120.00n L=30.00n
MM12 net3 net23 net040 VSS nch_mac W=120.00n L=30.00n
MM9 net7 net11 net044 VSS nch_mac W=120.00n L=30.00n
MM8 net23 net11 net7 VSS nch_mac W=120.00n L=30.00n
MM0 Z net19 VSS VSS nch_mac W=400.00n L=30.00n
MM5 net11 I VSS VSS nch_mac W=120.00n L=30.00n
MM14 net0103 net23 net083 VDD pch_mac W=200.00n L=30.00n
MM15 net083 net23 VDD VDD pch_mac W=200.00n L=30.00n
MM1 net087 net11 VDD VDD pch_mac W=200.00n L=30.00n
MM2 net0107 net11 net087 VDD pch_mac W=200.00n L=30.00n
MM11 net19 net23 net38 VDD pch_mac W=200.00n L=30.00n
MM10 net38 net23 net0103 VDD pch_mac W=200.00n L=30.00n
MM7 net42 net11 net0107 VDD pch_mac W=200.00n L=30.00n
MM6 net23 net11 net42 VDD pch_mac W=200.00n L=30.00n
MM3 Z net19 VDD VDD pch_mac W=400.00n L=30.00n
MM4 net11 I VDD VDD pch_mac W=200.00n L=30.00n
.ENDS DEL4V4
.SUBCKT DGRNQNV4 CK D QN RN VDD VSS
MM0 net156 c net163 VDD pch_mac W=200.00n L=30.00n
MM5 net152 net163 VDD VDD pch_mac W=200.00n L=30.00n
MM7 net163 cn net91 VDD pch_mac W=120.00n L=30.00n
MM8 net91 net152 VDD VDD pch_mac W=120.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM15 net152 cn net167 VDD pch_mac W=200.00n L=30.00n
MM19 net119 net128 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net167 c net119 VDD pch_mac W=120.00n L=30.00n
MM26 net156 RN VDD VDD pch_mac W=120.00n L=30.00n
MM27 net156 D VDD VDD pch_mac W=200.00n L=30.00n
MM21 net128 net167 VDD VDD pch_mac W=120.00n L=30.00n
MM23 QN net167 VDD VDD pch_mac W=400.00n L=30.00n
MM16 net144 net128 VSS VSS nch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM14 net152 c net167 VSS nch_mac W=200.00n L=30.00n
MM9 net136 net152 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net167 cn net144 VSS nch_mac W=120.00n L=30.00n
MM25 net156 D net148 VSS nch_mac W=200.00n L=30.00n
MM18 net128 net167 VSS VSS nch_mac W=120.00n L=30.00n
MM22 QN net167 VSS VSS nch_mac W=400.00n L=30.00n
MM6 net163 c net136 VSS nch_mac W=120.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM3 net156 cn net163 VSS nch_mac W=200.00n L=30.00n
MM24 net148 RN VSS VSS nch_mac W=200.00n L=30.00n
MM4 net152 net163 VSS VSS nch_mac W=200.00n L=30.00n
.ENDS DGRNQNV4
.SUBCKT DGRSNQNV4 CK D QN RN SN VDD VSS
MM28 net112 snn VDD VDD pch_mac W=200.00n L=30.00n
MM27 snn SN VDD VDD pch_mac W=120.00n L=30.00n
MM20 net188 c net100 VDD pch_mac W=120.00n L=30.00n
MM19 net100 net141 VDD VDD pch_mac W=120.00n L=30.00n
MM15 net169 cn net188 VDD pch_mac W=200.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM8 net136 net169 VDD VDD pch_mac W=120.00n L=30.00n
MM7 net192 cn net136 VDD pch_mac W=120.00n L=30.00n
MM5 net169 net192 VDD VDD pch_mac W=200.00n L=30.00n
MM0 net181 c net192 VDD pch_mac W=200.00n L=30.00n
MM23 QN net188 VDD VDD pch_mac W=400.00n L=30.00n
MM21 net141 net188 VDD VDD pch_mac W=120.00n L=30.00n
MM24 net181 RN VDD VDD pch_mac W=120.00n L=30.00n
MM1 net181 D net112 VDD pch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM26 snn SN VSS VSS nch_mac W=120.00n L=30.00n
MM16 net165 net141 VSS VSS nch_mac W=120.00n L=30.00n
MM29 net181 snn net177 VSS nch_mac W=120.00n L=30.00n
MM6 net192 c net173 VSS nch_mac W=120.00n L=30.00n
MM22 QN net188 VSS VSS nch_mac W=400.00n L=30.00n
MM18 net141 net188 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net188 cn net165 VSS nch_mac W=120.00n L=30.00n
MM14 net169 c net188 VSS nch_mac W=200.00n L=30.00n
MM25 net181 D net177 VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM3 net181 cn net192 VSS nch_mac W=200.00n L=30.00n
MM9 net173 net169 VSS VSS nch_mac W=120.00n L=30.00n
MM4 net169 net192 VSS VSS nch_mac W=200.00n L=30.00n
MM2 net177 RN VSS VSS nch_mac W=200.00n L=30.00n
.ENDS DGRSNQNV4
.SUBCKT DQNV4 CK D QN VDD VSS
MM14 net186 c net181 VSS nch_mac W=0.2u L=30.00n
MM3 net182 cn net177 VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM22 QN net181 VSS VSS nch_mac W=0.4u L=30.00n
MM16 net170 net190 VSS VSS nch_mac W=0.2u L=30.00n
MM2 net182 D VSS VSS nch_mac W=200.00n L=30.00n
MM4 net186 net177 VSS VSS nch_mac W=0.2u L=30.00n
MM18 net190 net181 VSS VSS nch_mac W=120.00n L=30.00n
MM9 net166 net186 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net181 cn net170 VSS nch_mac W=0.2u L=30.00n
MM6 net177 c net166 VSS nch_mac W=120.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM7 net177 cn net121 VDD pch_mac W=120.00n L=30.00n
MM19 net125 net190 VDD VDD pch_mac W=0.2u L=30.00n
MM8 net121 net186 VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM23 QN net181 VDD VDD pch_mac W=0.4u L=30.00n
MM21 net190 net181 VDD VDD pch_mac W=120.00n L=30.00n
MM5 net186 net177 VDD VDD pch_mac W=0.2u L=30.00n
MM1 net182 D VDD VDD pch_mac W=200.00n L=30.00n
MM15 net186 cn net181 VDD pch_mac W=0.2u L=30.00n
MM0 net182 c net177 VDD pch_mac W=0.2u L=30.00n
MM20 net181 c net125 VDD pch_mac W=0.2u L=30.00n
.ENDS DQNV4
.SUBCKT DQV4 CK D Q VDD VSS
MM24 net175 cn net191 VSS nch_mac W=120.00n L=30.00n
MM27 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM4 net156 cn net155 VSS nch_mac W=0.2u L=30.00n
MM0 net148 net155 VSS VSS nch_mac W=200.00n L=30.00n
MM11 VSS net148 net163 VSS nch_mac W=120.00n L=30.00n
MM17 s net191 VSS VSS nch_mac W=0.2u L=30.00n
MM30 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM5 net156 D VSS VSS nch_mac W=200.00n L=30.00n
MM12 net163 c net155 VSS nch_mac W=120.00n L=30.00n
MM3 net148 c net191 VSS nch_mac W=0.2u L=30.00n
MM42 Q s VSS VSS nch_mac W=0.4u L=30.00n
MM23 VSS s net175 VSS nch_mac W=120.00n L=30.00n
MM2 net148 cn net191 VDD pch_mac W=0.2u L=30.00n
MM25 net124 c net191 VDD pch_mac W=120.00n L=30.00n
MM7 net156 D VDD VDD pch_mac W=0.2u L=30.00n
MM1 net148 net155 VDD VDD pch_mac W=0.2u L=30.00n
MM13 VDD net148 net116 VDD pch_mac W=120.00n L=30.00n
MM18 s net191 VDD VDD pch_mac W=200.00n L=30.00n
MM43 Q s VDD VDD pch_mac W=0.4u L=30.00n
MM14 net116 cn net155 VDD pch_mac W=120.00n L=30.00n
MM6 net156 c net155 VDD pch_mac W=0.2u L=30.00n
MM28 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM26 VDD s net124 VDD pch_mac W=120.00n L=30.00n
MM29 c cn VDD VDD pch_mac W=0.2u L=30.00n
.ENDS DQV4
.SUBCKT DRNQNV4 CK D QN RDN VDD VSS
MM21 net150 net169 VDD VDD pch_mac W=200.00n L=30.00n
MM23 QN net170 VDD VDD pch_mac W=400.00n L=30.00n
MM19 net170 net150 VDD VDD pch_mac W=200.00n L=30.00n
MM20 net170 c net169 VDD pch_mac W=120.00n L=30.00n
MM15 net154 cn net169 VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM5 net154 net137 VDD VDD pch_mac W=0.2u L=30.00n
MM1 net142 D VDD VDD pch_mac W=0.2u L=30.00n
MM0 net142 c net137 VDD pch_mac W=0.2u L=30.00n
MM7 net137 cn net82 VDD pch_mac W=0.2u L=30.00n
MM8 net82 net154 VDD VDD pch_mac W=120.00n L=30.00n
MM25 net82 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM27 net150 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM24 net162 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM4 net154 net137 VSS VSS nch_mac W=0.2u L=30.00n
MM18 net150 RDN net146 VSS nch_mac W=200.00n L=30.00n
MM30 net146 net169 VSS VSS nch_mac W=200.00n L=30.00n
MM2 net142 D VSS VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM3 net142 cn net137 VSS nch_mac W=0.12u L=30.00n
MM9 net130 net154 net162 VSS nch_mac W=120.00n L=30.00n
MM6 net137 c net130 VSS nch_mac W=120.00n L=30.00n
MM22 QN net170 VSS VSS nch_mac W=400.00n L=30.00n
MM16 net170 net150 VSS VSS nch_mac W=200.00n L=30.00n
MM17 net170 cn net169 VSS nch_mac W=120.00n L=30.00n
MM14 net154 c net169 VSS nch_mac W=0.2u L=30.00n
.ENDS DRNQNV4
.SUBCKT DRNQV4 CK D Q RDN VDD VSS
MM14 net100 c net91 VSS nch_mac W=0.2u L=30.00n
MM17 net91 cn net80 VSS nch_mac W=120.00n L=30.00n
MM16 net80 net82 VSS VSS nch_mac W=120.00n L=30.00n
MM18 net82 RDN net72 VSS nch_mac W=0.2u L=30.00n
MM30 net72 net91 VSS VSS nch_mac W=0.2u L=30.00n
MM24 net92 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM6 net115 c net116 VSS nch_mac W=120.00n L=30.00n
MM22 Q net82 VSS VSS nch_mac W=0.4u L=30.00n
MM3 net104 cn net115 VSS nch_mac W=0.12u L=30.00n
MM9 net116 net100 net92 VSS nch_mac W=120.00n L=30.00n
MM2 net104 D VSS VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM4 net100 net115 VSS VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM23 Q net82 VDD VDD pch_mac W=0.4u L=30.00n
MM20 net91 c net143 VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM15 net100 cn net91 VDD pch_mac W=0.2u L=30.00n
MM19 net143 net82 VDD VDD pch_mac W=120.00n L=30.00n
MM1 net104 D VDD VDD pch_mac W=0.2u L=30.00n
MM7 net115 cn net128 VDD pch_mac W=0.2u L=30.00n
MM27 net82 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM25 net128 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM0 net104 c net115 VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM5 net100 net115 VDD VDD pch_mac W=0.2u L=30.00n
MM21 net82 net91 VDD VDD pch_mac W=0.2u L=30.00n
MM8 net128 net100 VDD VDD pch_mac W=120.00n L=30.00n
.ENDS DRNQV4
.SUBCKT DRQNV4 CK D QN RD VDD VSS
MM7 net144 cn net84 VDD pch_mac W=120.00n L=30.00n
MM1 net145 D VDD VDD pch_mac W=200.00n L=30.00n
MM15 net129 cn net136 VDD pch_mac W=200.00n L=30.00n
MM23 QN net136 VDD VDD pch_mac W=400.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM0 net145 c net144 VDD pch_mac W=200.00n L=30.00n
MM26 net88 RD VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM8 net84 net129 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net136 c net104 VDD pch_mac W=120.00n L=30.00n
MM24 net92 RD VDD VDD pch_mac W=200.00n L=30.00n
MM21 net179 net136 VDD VDD pch_mac W=120.00n L=30.00n
MM5 net129 net144 net92 VDD pch_mac W=200.00n L=30.00n
MM19 net104 net179 net88 VDD pch_mac W=120.00n L=30.00n
MM27 net136 RD VSS VSS nch_mac W=120.00n L=30.00n
MM22 QN net136 VSS VSS nch_mac W=400.00n L=30.00n
MM3 net145 cn net144 VSS nch_mac W=200.00n L=30.00n
MM9 net137 net129 VSS VSS nch_mac W=120.00n L=30.00n
MM18 net179 net136 VSS VSS nch_mac W=120.00n L=30.00n
MM25 net129 RD VSS VSS nch_mac W=120.00n L=30.00n
MM2 net145 D VSS VSS nch_mac W=200.00n L=30.00n
MM14 net129 c net136 VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM4 net129 net144 VSS VSS nch_mac W=200.00n L=30.00n
MM17 net136 cn net177 VSS nch_mac W=120.00n L=30.00n
MM16 net177 net179 VSS VSS nch_mac W=120.00n L=30.00n
MM6 net144 c net137 VSS nch_mac W=120.00n L=30.00n
.ENDS DRQNV4
.SUBCKT DRQV4 CK D Q RD VDD VSS
MM16 net185 net187 VSS VSS nch_mac W=120.00n L=30.00n
MM28 Q net187 VSS VSS nch_mac W=400.00n L=30.00n
MM6 net192 c net177 VSS nch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM27 net196 RD VSS VSS nch_mac W=120.00n L=30.00n
MM18 net187 net196 VSS VSS nch_mac W=200.00n L=30.00n
MM25 net201 RD VSS VSS nch_mac W=120.00n L=30.00n
MM2 net197 D VSS VSS nch_mac W=200.00n L=30.00n
MM3 net197 cn net192 VSS nch_mac W=200.00n L=30.00n
MM9 net177 net201 VSS VSS nch_mac W=120.00n L=30.00n
MM14 net201 c net196 VSS nch_mac W=200.00n L=30.00n
MM4 net201 net192 VSS VSS nch_mac W=200.00n L=30.00n
MM17 net196 cn net185 VSS nch_mac W=120.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM29 Q net187 VDD VDD pch_mac W=400.00n L=30.00n
MM0 net197 c net192 VDD pch_mac W=200.00n L=30.00n
MM26 net128 RD VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM8 net124 net201 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net196 c net132 VDD pch_mac W=120.00n L=30.00n
MM24 net152 RD VDD VDD pch_mac W=200.00n L=30.00n
MM21 net187 net196 VDD VDD pch_mac W=200.00n L=30.00n
MM5 net201 net192 net152 VDD pch_mac W=200.00n L=30.00n
MM19 net132 net187 net128 VDD pch_mac W=120.00n L=30.00n
MM7 net192 cn net124 VDD pch_mac W=120.00n L=30.00n
MM1 net197 D VDD VDD pch_mac W=200.00n L=30.00n
MM15 net201 cn net196 VDD pch_mac W=200.00n L=30.00n
.ENDS DRQV4
.SUBCKT DSRNQV4 CK D Q RDN SDN VDD VSS
MM15 net170 cn net181 VDD pch_mac W=200.00n L=30.00n
MM23 Q net146 VDD VDD pch_mac W=400.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM19 net130 net146 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net181 c net130 VDD pch_mac W=120.00n L=30.00n
MM24 net170 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM5 net170 net185 VDD VDD pch_mac W=200.00n L=30.00n
MM21 net146 net181 VDD VDD pch_mac W=200.00n L=30.00n
MM8 net185 cn net86 VDD pch_mac W=120.00n L=30.00n
MM37 net130 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM35 net86 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM1 net174 D VDD VDD pch_mac W=120.00n L=30.00n
MM36 net86 net170 VDD VDD pch_mac W=120.00n L=30.00n
MM27 net146 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM0 net174 c net185 VDD pch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM17 net181 cn net198 VSS nch_mac W=120.00n L=30.00n
MM4 net170 net185 net162 VSS nch_mac W=200.00n L=30.00n
MM16 net198 net146 net186 VSS nch_mac W=120.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM29 net186 SDN VSS VSS nch_mac W=120.00n L=30.00n
MM3 net174 cn net185 VSS nch_mac W=120.00n L=30.00n
MM14 net170 c net181 VSS nch_mac W=200.00n L=30.00n
MM2 net174 D VSS VSS nch_mac W=120.00n L=30.00n
MM22 Q net146 VSS VSS nch_mac W=400.00n L=30.00n
MM26 net162 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM6 net158 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM7 net185 c net150 VSS nch_mac W=120.00n L=30.00n
MM9 net150 net170 net158 VSS nch_mac W=120.00n L=30.00n
MM18 net146 RDN net142 VSS nch_mac W=200.00n L=30.00n
MM30 net142 net181 VSS VSS nch_mac W=200.00n L=30.00n
.ENDS DSRNQV4
.SUBCKT DSNQNV4 CK D QN SDN VDD VSS
MM21 net161 net156 VDD VDD pch_mac W=120.00n L=30.00n
MM19 net117 net161 VDD VDD pch_mac W=0.2u L=30.00n
MM1 net125 D VDD VDD pch_mac W=0.2u L=30.00n
MM20 net156 c net117 VDD pch_mac W=0.2u L=30.00n
MM5 net133 net132 VDD VDD pch_mac W=0.2u L=30.00n
MM0 net125 c net132 VDD pch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM23 QN net156 VDD VDD pch_mac W=0.4u L=30.00n
MM29 net117 SDN VDD VDD pch_mac W=0.2u L=30.00n
MM7 net132 cn net84 VDD pch_mac W=120.00n L=30.00n
MM8 net84 net133 VDD VDD pch_mac W=120.00n L=30.00n
MM28 net133 SDN VDD VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM15 net133 cn net156 VDD pch_mac W=0.2u L=30.00n
MM25 net165 net161 VSS VSS nch_mac W=0.2u L=30.00n
MM22 QN net156 VSS VSS nch_mac W=0.4u L=30.00n
MM18 net161 net156 VSS VSS nch_mac W=120.00n L=30.00n
MM2 net125 D VSS VSS nch_mac W=0.2u L=30.00n
MM3 net125 cn net132 VSS nch_mac W=0.2u L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM17 net156 cn net169 VSS nch_mac W=0.2u L=30.00n
MM16 net169 SDN net165 VSS nch_mac W=0.2u L=30.00n
MM9 net141 net133 VSS VSS nch_mac W=120.00n L=30.00n
MM4 net133 net132 net157 VSS nch_mac W=200.00n L=30.00n
MM24 net157 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM14 net133 c net156 VSS nch_mac W=0.2u L=30.00n
MM6 net132 c net141 VSS nch_mac W=120.00n L=30.00n
.ENDS DSNQNV4
.SUBCKT DSNQV4 CK D Q SDN VDD VSS
MM17 net208 cn net189 VSS nch_mac W=120.00n L=30.00n
MM16 net189 net197 net193 VSS nch_mac W=120.00n L=30.00n
MM14 net225 c net208 VSS nch_mac W=0.2u L=30.00n
MM22 Q net197 VSS VSS nch_mac W=0.4u L=30.00n
MM25 net193 SDN VSS VSS nch_mac W=120.00n L=30.00n
MM3 net233 cn net232 VSS nch_mac W=0.2u L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM4 net225 net232 net201 VSS nch_mac W=200.00n L=30.00n
MM9 net217 net225 VSS VSS nch_mac W=120.00n L=30.00n
MM6 net232 c net217 VSS nch_mac W=120.00n L=30.00n
MM18 net197 net208 VSS VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM24 net201 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM2 net233 D VSS VSS nch_mac W=0.2u L=30.00n
MM8 net140 net225 VDD VDD pch_mac W=120.00n L=30.00n
MM21 net197 net208 VDD VDD pch_mac W=0.2u L=30.00n
MM19 net241 net197 VDD VDD pch_mac W=120.00n L=30.00n
MM28 net225 SDN VDD VDD pch_mac W=0.2u L=30.00n
MM23 Q net197 VDD VDD pch_mac W=0.4u L=30.00n
MM29 net241 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM1 net233 D VDD VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM7 net232 cn net140 VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM20 net208 c net241 VDD pch_mac W=120.00n L=30.00n
MM15 net225 cn net208 VDD pch_mac W=0.2u L=30.00n
MM5 net225 net232 VDD VDD pch_mac W=0.2u L=30.00n
MM0 net233 c net232 VDD pch_mac W=0.2u L=30.00n
.ENDS DSNQV4
.SUBCKT EDRNQNV4 CK D E QN RDN VDD VSS
MM7 net198 cn net98 VDD pch_mac W=120.00n L=30.00n
MM21 net193 s VDD VDD pch_mac W=120.00n L=30.00n
MM5 net215 net198 net90 VDD pch_mac W=200.00n L=30.00n
MM15 net215 cn s VDD pch_mac W=200.00n L=30.00n
MM23 QN s VDD VDD pch_mac W=400.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM34 net138 en VDD VDD pch_mac W=200.00n L=30.00n
MM35 net223 E net146 VDD pch_mac W=120.00n L=30.00n
MM36 net146 s VDD VDD pch_mac W=120.00n L=30.00n
MM37 net223 D net138 VDD pch_mac W=200.00n L=30.00n
MM39 en E VDD VDD pch_mac W=120.00n L=30.00n
MM0 net223 c net198 VDD pch_mac W=200.00n L=30.00n
MM26 net106 R VDD VDD pch_mac W=120.00n L=30.00n
MM28 R RDN VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM8 net98 net215 VDD VDD pch_mac W=120.00n L=30.00n
MM20 s c net110 VDD pch_mac W=120.00n L=30.00n
MM19 net110 net193 net106 VDD pch_mac W=120.00n L=30.00n
MM24 net90 R VDD VDD pch_mac W=200.00n L=30.00n
MM25 net215 R VSS VSS nch_mac W=120.00n L=30.00n
MM3 net223 cn net198 VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM32 net223 en net187 VSS nch_mac W=120.00n L=30.00n
MM16 net191 net193 VSS VSS nch_mac W=120.00n L=30.00n
MM33 net187 s VSS VSS nch_mac W=120.00n L=30.00n
MM27 s R VSS VSS nch_mac W=120.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM38 en E VSS VSS nch_mac W=120.00n L=30.00n
MM31 net183 E VSS VSS nch_mac W=200.00n L=30.00n
MM29 R RDN VSS VSS nch_mac W=120.00n L=30.00n
MM22 QN s VSS VSS nch_mac W=400.00n L=30.00n
MM9 net231 net215 VSS VSS nch_mac W=120.00n L=30.00n
MM14 net215 c s VSS nch_mac W=200.00n L=30.00n
MM30 net223 D net183 VSS nch_mac W=200.00n L=30.00n
MM18 net193 s VSS VSS nch_mac W=120.00n L=30.00n
MM4 net215 net198 VSS VSS nch_mac W=200.00n L=30.00n
MM17 s cn net191 VSS nch_mac W=120.00n L=30.00n
MM6 net198 c net231 VSS nch_mac W=120.00n L=30.00n
.ENDS EDRNQNV4
.SUBCKT INV4 I ZN VDD VSS
MM2 ZN I VSS VSS nch_mac W=0.4u L=30.00n
MM3 ZN I VDD VDD pch_mac W=0.4u L=30.00n
.ENDS INV4
.SUBCKT LAHQV4 D E Q VDD VSS
MM12 net51 EN VDD VDD pch_mac W=200.00n L=30.00n
MM3 ENN EN VDD VDD pch_mac W=0.2u L=30.00n
MM8 net59 net72 VDD VDD pch_mac W=120.00n L=30.00n
MM7 net80 ENN net59 VDD pch_mac W=120.00n L=30.00n
MM14 Q net80 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net80 D net51 VDD pch_mac W=200.00n L=30.00n
MM11 EN E VDD VDD pch_mac W=120.00n L=30.00n
MM5 net72 net80 VDD VDD pch_mac W=120.00n L=30.00n
MM10 EN E VSS VSS nch_mac W=120.00n L=30.00n
MM9 net92 EN VSS VSS nch_mac W=120.00n L=30.00n
MM6 net80 net72 net92 VSS nch_mac W=120.00n L=30.00n
MM13 net100 D VSS VSS nch_mac W=200.00n L=30.00n
MM2 net80 ENN net100 VSS nch_mac W=0.2u L=30.00n
MM4 net72 net80 VSS VSS nch_mac W=120.00n L=30.00n
MM0 ENN EN VSS VSS nch_mac W=0.2u L=30.00n
MM15 Q net80 VSS VSS nch_mac W=0.4u L=30.00n
.ENDS LAHQV4
.SUBCKT LAHRNQV4 D E Q RDN VDD VSS
MM1 net67 EN VDD VDD pch_mac W=200.00n L=30.00n
MM12 net108 D net67 VDD pch_mac W=200.00n L=30.00n
MM19 net108 RDN VDD VDD pch_mac W=200.00n L=30.00n
MM5 net92 net108 VDD VDD pch_mac W=120.00n L=30.00n
MM8 net51 net92 VDD VDD pch_mac W=120.00n L=30.00n
MM7 net108 ENN net51 VDD pch_mac W=120.00n L=30.00n
MM14 Q net108 VDD VDD pch_mac W=0.4u L=30.00n
MM3 ENN EN VDD VDD pch_mac W=0.2u L=30.00n
MM11 EN E VDD VDD pch_mac W=120.00n L=30.00n
MM15 Q net108 VSS VSS nch_mac W=0.4u L=30.00n
MM0 ENN EN VSS VSS nch_mac W=0.2u L=30.00n
MM16 net104 RDN VSS VSS nch_mac W=200.00n L=30.00n
MM10 EN E VSS VSS nch_mac W=120.00n L=30.00n
MM2 net100 D net104 VSS nch_mac W=200.00n L=30.00n
MM4 net92 net108 VSS VSS nch_mac W=120.00n L=30.00n
MM18 net96 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM9 net88 EN net96 VSS nch_mac W=120.00n L=30.00n
MM13 net108 ENN net100 VSS nch_mac W=0.2u L=30.00n
MM6 net108 net92 net88 VSS nch_mac W=120.00n L=30.00n
.ENDS LAHRNQV4
.SUBCKT LAHRSNQV4 D E Q RDN SDN VDD VSS
MM23 Q pm VDD VDD pch_mac W=400.00n L=30.00n
MM14 net114 D net106 VDD pch_mac W=120.00n L=30.00n
MM26 pm E net98 VDD pch_mac W=120.00n L=30.00n
MM20 EN E VDD VDD pch_mac W=120.00n L=30.00n
MM18 net147 pm VDD VDD pch_mac W=120.00n L=30.00n
MM17 pm s net118 VDD pch_mac W=120.00n L=30.00n
MM15 pm EN net114 VDD pch_mac W=120.00n L=30.00n
MM16 net118 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM24 net94 net147 VDD VDD pch_mac W=120.00n L=30.00n
MM25 net98 s net94 VDD pch_mac W=120.00n L=30.00n
MM22 s SDN VDD VDD pch_mac W=120.00n L=30.00n
MM13 net106 s VDD VDD pch_mac W=120.00n L=30.00n
MM9 net147 pm VSS VSS nch_mac W=120.00n L=30.00n
MM7 pm E net159 VSS nch_mac W=120.00n L=30.00n
MM8 pm s VSS VSS nch_mac W=120.00n L=30.00n
MM6 net159 D net163 VSS nch_mac W=120.00n L=30.00n
MM5 net163 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM1 Q pm VSS VSS nch_mac W=400.00n L=30.00n
MM4 EN E VSS VSS nch_mac W=120.00n L=30.00n
MM2 s SDN VSS VSS nch_mac W=120.00n L=30.00n
MM11 net139 net147 net143 VSS nch_mac W=120.00n L=30.00n
MM10 net143 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM12 pm EN net139 VSS nch_mac W=120.00n L=30.00n
.ENDS LAHRSNQV4
.SUBCKT LAHSQV4 D E Q SD VDD VSS
MM17 ENN EN VDD VDD pch_mac W=0.2u L=30.00n
MM11 EN E VDD VDD pch_mac W=0.12u L=30.00n
MM14 Q net169 VDD VDD pch_mac W=0.4u L=30.00n
MM19 net136 SD VDD VDD pch_mac W=200.00n L=30.00n
MM18 net132 EN net136 VDD pch_mac W=200.00n L=30.00n
MM1 net169 D net132 VDD pch_mac W=200.00n L=30.00n
MM5 net165 net169 VDD VDD pch_mac W=0.12u L=30.00n
MM21 net156 SD VDD VDD pch_mac W=120.00n L=30.00n
MM7 net169 ENN net160 VDD pch_mac W=120.00n L=30.00n
MM8 net160 net165 net156 VDD pch_mac W=120.00n L=30.00n
MM10 EN E VSS VSS nch_mac W=0.12u L=30.00n
MM2 net169 ENN net173 VSS nch_mac W=0.2u L=30.00n
MM9 net193 EN VSS VSS nch_mac W=120.00n L=30.00n
MM6 net169 net165 net193 VSS nch_mac W=120.00n L=30.00n
MM20 net173 D VSS VSS nch_mac W=0.2u L=30.00n
MM13 ENN EN VSS VSS nch_mac W=0.2u L=30.00n
MM22 net169 SD VSS VSS nch_mac W=0.12u L=30.00n
MM15 Q net169 VSS VSS nch_mac W=0.4u L=30.00n
MM4 net165 net169 VSS VSS nch_mac W=0.12u L=30.00n
.ENDS LAHSQV4
.SUBCKT LALQV4 D EN Q VDD VSS
MM23 Q net88 VDD VDD pch_mac W=0.4u L=30.00n
MM11 ENN EN VDD VDD pch_mac W=0.12u L=30.00n
MM13 ENNN ENN VDD VDD pch_mac W=0.2u L=30.00n
MM1 net88 ENNN net59 VDD pch_mac W=0.2u L=30.00n
MM14 net59 D VDD VDD pch_mac W=0.2u L=30.00n
MM7 net88 net76 net67 VDD pch_mac W=120.00n L=30.00n
MM8 net67 ENN VDD VDD pch_mac W=120.00n L=30.00n
MM5 net76 net88 VDD VDD pch_mac W=120.00n L=30.00n
MM4 net76 net88 VSS VSS nch_mac W=120.00n L=30.00n
MM22 Q net88 VSS VSS nch_mac W=0.4u L=30.00n
MM12 ENNN ENN VSS VSS nch_mac W=0.2u L=30.00n
MM6 net88 ENNN net100 VSS nch_mac W=120.00n L=30.00n
MM15 net92 ENN VSS VSS nch_mac W=0.2u L=30.00n
MM2 net88 D net92 VSS nch_mac W=0.2u L=30.00n
MM9 net100 net76 VSS VSS nch_mac W=120.00n L=30.00n
MM10 ENN EN VSS VSS nch_mac W=120.00n L=30.00n
.ENDS LALQV4
.SUBCKT LALRNQV4 D EN Q RDN VDD VSS
MM11 ENN EN VDD VDD pch_mac W=120.00n L=30.00n
MM17 net102 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM12 net102 D net69 VDD pch_mac W=200.00n L=30.00n
MM1 net69 EN VDD VDD pch_mac W=200.00n L=30.00n
MM7 net102 ENN net61 VDD pch_mac W=120.00n L=30.00n
MM14 Q net102 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net90 net102 VDD VDD pch_mac W=120.00n L=30.00n
MM8 net61 net90 VDD VDD pch_mac W=120.00n L=30.00n
MM10 ENN EN VSS VSS nch_mac W=120.00n L=30.00n
MM4 net90 net102 VSS VSS nch_mac W=120.00n L=30.00n
MM9 net86 EN net94 VSS nch_mac W=120.00n L=30.00n
MM6 net102 net90 net86 VSS nch_mac W=120.00n L=30.00n
MM15 Q net102 VSS VSS nch_mac W=400.00n L=30.00n
MM2 net98 D net106 VSS nch_mac W=200.00n L=30.00n
MM18 net94 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM16 net106 RDN VSS VSS nch_mac W=200.00n L=30.00n
MM13 net102 ENN net98 VSS nch_mac W=200.00n L=30.00n
.ENDS LALRNQV4
.SUBCKT LALRSNQV4 D EN Q RDN SDN VDD VSS
MM15 pm EN net106 VDD pch_mac W=120.00n L=30.00n
MM16 net98 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM17 pm s net98 VDD pch_mac W=120.00n L=30.00n
MM22 s SDN VDD VDD pch_mac W=120.00n L=30.00n
MM23 Q pm VDD VDD pch_mac W=400.00n L=30.00n
MM18 net167 pm VDD VDD pch_mac W=120.00n L=30.00n
MM20 ENN EN VDD VDD pch_mac W=120.00n L=30.00n
MM24 net122 net167 VDD VDD pch_mac W=120.00n L=30.00n
MM25 net118 s net122 VDD pch_mac W=120.00n L=30.00n
MM26 pm ENN net118 VDD pch_mac W=120.00n L=30.00n
MM13 net110 s VDD VDD pch_mac W=120.00n L=30.00n
MM14 net106 D net110 VDD pch_mac W=120.00n L=30.00n
MM4 ENN EN VSS VSS nch_mac W=120.00n L=30.00n
MM5 net139 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM6 net135 D net139 VSS nch_mac W=120.00n L=30.00n
MM7 pm ENN net135 VSS nch_mac W=120.00n L=30.00n
MM8 pm s VSS VSS nch_mac W=120.00n L=30.00n
MM9 net167 pm VSS VSS nch_mac W=120.00n L=30.00n
MM10 net163 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM11 net159 net167 net163 VSS nch_mac W=120.00n L=30.00n
MM12 pm EN net159 VSS nch_mac W=120.00n L=30.00n
MM1 Q pm VSS VSS nch_mac W=400.00n L=30.00n
MM2 s SDN VSS VSS nch_mac W=120.00n L=30.00n
.ENDS LALRSNQV4
.SUBCKT LALSNQV4 D EN Q SDN VDD VSS
MM18 S SDN VDD VDD pch_mac W=0.12u L=30.00n
MM11 ENN EN VDD VDD pch_mac W=0.12u L=30.00n
MM21 net112 ENNN net79 VDD pch_mac W=200.00n L=30.00n
MM12 net71 S VDD VDD pch_mac W=200.00n L=30.00n
MM1 net79 D net71 VDD pch_mac W=200.00n L=30.00n
MM14 Q net112 VDD VDD pch_mac W=0.4u L=30.00n
MM7 net112 net104 net63 VDD pch_mac W=120.00n L=30.00n
MM8 net63 ENN net59 VDD pch_mac W=120.00n L=30.00n
MM13 net59 S VDD VDD pch_mac W=120.00n L=30.00n
MM5 net104 net112 VDD VDD pch_mac W=120.00n L=30.00n
MM20 ENNN ENN VDD VDD pch_mac W=0.2u L=30.00n
MM17 S SDN VSS VSS nch_mac W=120.00n L=30.00n
MM19 ENNN ENN VSS VSS nch_mac W=0.2u L=30.00n
MM10 ENN EN VSS VSS nch_mac W=120.00n L=30.00n
MM22 net112 S VSS VSS nch_mac W=200.00n L=30.00n
MM2 net112 D net116 VSS nch_mac W=200.00n L=30.00n
MM9 net92 net104 VSS VSS nch_mac W=120.00n L=30.00n
MM6 net112 ENNN net92 VSS nch_mac W=120.00n L=30.00n
MM4 net104 net112 VSS VSS nch_mac W=120.00n L=30.00n
MM23 net116 ENN VSS VSS nch_mac W=200.00n L=30.00n
MM15 Q net112 VSS VSS nch_mac W=0.4u L=30.00n
.ENDS LALSNQV4
.SUBCKT MAJ23V4 A1 A2 A3 Z VDD VSS
MM9 net13 A2 VSS VSS nch_mac W=200.00n L=30.00n
MM8 net21 A1 net13 VSS nch_mac W=200.00n L=30.00n
MM5 net9 A2 VSS VSS nch_mac W=200.00n L=30.00n
MM2 net9 A1 VSS VSS nch_mac W=200.00n L=30.00n
MM4 net21 A3 net9 VSS nch_mac W=200.00n L=30.00n
MM11 Z net21 VSS VSS nch_mac W=400.00n L=30.00n
MM10 Z net21 VDD VDD pch_mac W=400.00n L=30.00n
MM7 net21 A1 net32 VDD pch_mac W=200.00n L=30.00n
MM6 net32 A2 VDD VDD pch_mac W=200.00n L=30.00n
MM3 net21 A3 net49 VDD pch_mac W=200.00n L=30.00n
MM0 net49 A2 VDD VDD pch_mac W=200.00n L=30.00n
MM1 net49 A1 VDD VDD pch_mac W=200.00n L=30.00n
.ENDS MAJ23V4
.SUBCKT MUX2NV4 I0 I1 S ZN VDD VSS
MM36 net39 net43 ZN VSS nch_mac W=400.00n L=30.00n
MM47 net41 S ZN VSS nch_mac W=400.00n L=30.00n
MM49 net39 I0 VSS VSS nch_mac W=400.00n L=30.00n
MM31 net41 I1 VSS VSS nch_mac W=400.00n L=30.00n
MM53 net43 S VSS VSS nch_mac W=120.00n L=30.00n
MM54 net43 S VDD VDD pch_mac W=120.00n L=30.00n
MM39 net39 S ZN VDD pch_mac W=400.00n L=30.00n
MM50 net39 I0 VDD VDD pch_mac W=400.00n L=30.00n
MM32 net41 I1 VDD VDD pch_mac W=400.00n L=30.00n
MM48 net41 net43 ZN VDD pch_mac W=400.00n L=30.00n
.ENDS MUX2NV4
.SUBCKT MUX2V4 I0 I1 S Z VDD VSS
MM31 net41 I1 VSS VSS nch_mac W=160.00n L=30.00n
MM49 net39 I0 VSS VSS nch_mac W=160.00n L=30.00n
MM51 Z net_65 VSS VSS nch_mac W=400.00n L=30.00n
MM47 net41 S net_65 VSS nch_mac W=200.00n L=30.00n
MM36 net39 net43 net_65 VSS nch_mac W=160.00n L=30.00n
MM53 net43 S VSS VSS nch_mac W=120.00n L=30.00n
MM39 net39 S net_65 VDD pch_mac W=160.00n L=30.00n
MM54 net43 S VDD VDD pch_mac W=120.00n L=30.00n
MM32 net41 I1 VDD VDD pch_mac W=160.00n L=30.00n
MM48 net41 net43 net_65 VDD pch_mac W=160.00n L=30.00n
MM52 Z net_65 VDD VDD pch_mac W=400.00n L=30.00n
MM50 net39 I0 VDD VDD pch_mac W=160.00n L=30.00n
.ENDS MUX2V4
.SUBCKT MUX3NV4 I0 I1 I2 S0 S1 ZN VDD VSS
MM22 net114 net109 VSS VSS nch_mac W=200.00n L=30.00n
MM9 net90 S0N net109 VSS nch_mac W=200.00n L=30.00n
MM14 ZN net129 VSS VSS nch_mac W=400.00n L=30.00n
MM10 net94 S0 net109 VSS nch_mac W=200.00n L=30.00n
MM1 net98 I2 VSS VSS nch_mac W=200.00n L=30.00n
MM4 net94 I1 VSS VSS nch_mac W=200.00n L=30.00n
MM3 net90 I0 VSS VSS nch_mac W=120.00n L=30.00n
MM17 S0N S0 VSS VSS nch_mac W=120.00n L=30.00n
MM18 S1N S1 VSS VSS nch_mac W=120.00n L=30.00n
MM0 net122 S1 net129 VSS nch_mac W=200.00n L=30.00n
MM21 net122 net98 VSS VSS nch_mac W=200.00n L=30.00n
MM12 net114 S1N net129 VSS nch_mac W=200.00n L=30.00n
MM15 ZN net129 VDD VDD pch_mac W=400.00n L=30.00n
MM13 net114 S1 net129 VDD pch_mac W=200.00n L=30.00n
MM20 net122 net98 VDD VDD pch_mac W=200.00n L=30.00n
MM16 S0N S0 VDD VDD pch_mac W=120.00n L=30.00n
MM5 net94 I1 VDD VDD pch_mac W=200.00n L=30.00n
MM19 S1N S1 VDD VDD pch_mac W=120.00n L=30.00n
MM7 net98 I2 VDD VDD pch_mac W=200.00n L=30.00n
MM2 net90 I0 VDD VDD pch_mac W=120.00n L=30.00n
MM11 net94 S0N net109 VDD pch_mac W=200.00n L=30.00n
MM23 net114 net109 VDD VDD pch_mac W=200.00n L=30.00n
M200.00n net90 S0 net109 VDD pch_mac W=200.00n L=30.00n
MM6 net122 S1N net129 VDD pch_mac W=200.00n L=30.00n
.ENDS MUX3NV4
.SUBCKT MUX3V4 I0 I1 I2 S0 S1 Z VDD VSS
MM1 net100 I2 VSS VSS nch_mac W=200.00n L=30.00n
MM0 net100 S1 net95 VSS nch_mac W=200.00n L=30.00n
MM17 S0N S0 VSS VSS nch_mac W=120.00n L=30.00n
MM18 S1N S1 VSS VSS nch_mac W=120.00n L=30.00n
MM9 net80 S0N net107 VSS nch_mac W=200.00n L=30.00n
MM12 net107 S1N net95 VSS nch_mac W=200.00n L=30.00n
MM4 net76 I1 VSS VSS nch_mac W=200.00n L=30.00n
MM3 net80 I0 VSS VSS nch_mac W=120.00n L=30.00n
MM14 Z net95 VSS VSS nch_mac W=400.00n L=30.00n
MM10 net76 S0 net107 VSS nch_mac W=200.00n L=30.00n
MM19 S1N S1 VDD VDD pch_mac W=120.00n L=30.00n
MM6 net100 S1N net95 VDD pch_mac W=200.00n L=30.00n
MM13 net107 S1 net95 VDD pch_mac W=200.00n L=30.00n
MM2 net80 I0 VDD VDD pch_mac W=120.00n L=30.00n
MM16 S0N S0 VDD VDD pch_mac W=120.00n L=30.00n
MM8 net80 S0 net107 VDD pch_mac W=200.00n L=30.00n
MM15 Z net95 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net76 I1 VDD VDD pch_mac W=200.00n L=30.00n
MM7 net100 I2 VDD VDD pch_mac W=200.00n L=30.00n
MM11 net76 S0N net107 VDD pch_mac W=200.00n L=30.00n
.ENDS MUX3V4
.SUBCKT NAND2V4 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VSS nch_mac W=0.4u L=30.00n
MMN1 net18 A2 VSS VSS nch_mac W=0.4u L=30.00n
MM0 ZN A2 VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS NAND2V4
.SUBCKT NAND2XBV4 A1 B1 ZN VDD VSS
MM3 A1N A1 VSS VSS nch_mac W=0.175u L=30.00n
MM1 ZN B1 net18 VSS nch_mac W=0.4u L=30.00n
MMN1 net18 A1N VSS VSS nch_mac W=0.4u L=30.00n
MM4 A1N A1 VDD VDD pch_mac W=0.175u L=30.00n
MM0 ZN B1 VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1N VDD VDD pch_mac W=0.4u L=30.00n
.ENDS NAND2XBV4
.SUBCKT NAND3BBV4 A1 A2 B ZN VDD VSS
MM0 ZN A1N net028 VSS nch_mac W=0.4u L=30.00n
MM7 net028 A2N net9 VSS nch_mac W=0.4u L=30.00n
MM6 net9 B VSS VSS nch_mac W=0.4u L=30.00n
MM4 A1N A1 VSS VSS nch_mac W=0.175u L=30.00n
MM8 A2N A2 VSS VSS nch_mac W=0.175u L=30.00n
MM2 ZN A1N VDD VDD pch_mac W=0.38u L=30.00n
MM3 ZN A2N VDD VDD pch_mac W=0.38u L=30.00n
MM1 ZN B VDD VDD pch_mac W=0.4u L=30.00n
MM9 A2N A2 VDD VDD pch_mac W=0.175u L=30.00n
MM5 A1N A1 VDD VDD pch_mac W=0.175u L=30.00n
.ENDS NAND3BBV4
.SUBCKT NAND3V4 A1 A2 A3 ZN VDD VSS
MM1 ZN A1 net18 VSS nch_mac W=0.4u L=30.00n
MM3 net022 A3 VSS VSS nch_mac W=0.4u L=30.00n
MMN1 net18 A2 net022 VSS nch_mac W=0.4u L=30.00n
MM2 ZN A3 VDD VDD pch_mac W=0.4u L=30.00n
MM0 ZN A2 VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS NAND3V4
.SUBCKT NAND4BBV4 A1 A2 B1 B2 ZN VDD VSS
MM5 net92 B2 VSS VSS nch_mac W=400.00n L=30.00n
MM9 net76 A2 VSS VSS nch_mac W=200.00n L=30.00n
MM8 net76 A1 VSS VSS nch_mac W=200.00n L=30.00n
MM6 net88 B1 net92 VSS nch_mac W=400.00n L=30.00n
MM7 ZN net76 net88 VSS nch_mac W=400.00n L=30.00n
MM4 ZN net76 VDD VDD pch_mac W=400.00n L=30.00n
MM2 net76 A1 net63 VDD pch_mac W=200.00n L=30.00n
MM0 net63 A2 VDD VDD pch_mac W=200.00n L=30.00n
MM1 ZN B2 VDD VDD pch_mac W=400.00n L=30.00n
MM3 ZN B1 VDD VDD pch_mac W=400.00n L=30.00n
.ENDS NAND4BBV4
.SUBCKT NAND4V4 A1 A2 A3 A4 ZN VDD VSS
MM4 net026 A4 VSS VSS nch_mac W=0.39u L=30.00n
MM1 ZN A1 net18 VSS nch_mac W=0.39u L=30.00n
MM3 net022 A3 net026 VSS nch_mac W=0.39u L=30.00n
MMN1 net18 A2 net022 VSS nch_mac W=0.39u L=30.00n
MM5 ZN A4 VDD VDD pch_mac W=0.24u L=30.00n
MM2 ZN A3 VDD VDD pch_mac W=0.24u L=30.00n
MM0 ZN A2 VDD VDD pch_mac W=0.24u L=30.00n
MMP1 ZN A1 VDD VDD pch_mac W=0.24u L=30.00n
.ENDS NAND4V4
.SUBCKT NAND4XXBBV4 A1 A2 B1 B2 ZN VDD VSS
MM5 net92 net035 VSS VSS nch_mac W=0.4u L=30.00n
MM9 net035 A2 VSS VSS nch_mac W=0.175u L=30.00n
MM8 net035 A1 VSS VSS nch_mac W=0.175u L=30.00n
MM6 net88 B2 net92 VSS nch_mac W=0.4u L=30.00n
MM7 ZN B1 net88 VSS nch_mac W=0.4u L=30.00n
MM4 ZN net035 VDD VDD pch_mac W=0.4u L=30.00n
MM2 net035 A1 net63 VDD pch_mac W=0.175u L=30.00n
MM0 net63 A2 VDD VDD pch_mac W=0.175u L=30.00n
MM1 ZN B2 VDD VDD pch_mac W=0.4u L=30.00n
MM3 ZN B1 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS NAND4XXBBV4
.SUBCKT NDQV4 CKN D Q VDD VSS
MM2 net24 D VSS VSS nch_mac W=0.2u L=30.00n
MM3 net24 cn net35 VSS nch_mac W=0.2u L=30.00n
MM4 net20 net35 VSS VSS nch_mac W=0.2u L=30.00n
MM6 net35 c net40 VSS nch_mac W=120.00n L=30.00n
MM9 net40 net20 VSS VSS nch_mac W=120.00n L=30.00n
MM10 c CKN VSS VSS nch_mac W=0.2u L=30.00n
MM12 cn c VSS VSS nch_mac W=0.2u L=30.00n
MM14 net20 c net31 VSS nch_mac W=0.2u L=30.00n
MM16 net36 net16 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net31 cn net36 VSS nch_mac W=120.00n L=30.00n
MM18 net16 net31 VSS VSS nch_mac W=0.2u L=30.00n
MM22 Q net16 VSS VSS nch_mac W=0.4u L=30.00n
MM1 net24 D VDD VDD pch_mac W=0.2u L=30.00n
MM0 net24 c net35 VDD pch_mac W=0.2u L=30.00n
MM5 net20 net35 VDD VDD pch_mac W=0.2u L=30.00n
MM7 net35 cn net91 VDD pch_mac W=120.00n L=30.00n
MM8 net91 net20 VDD VDD pch_mac W=120.00n L=30.00n
MM11 c CKN VDD VDD pch_mac W=0.2u L=30.00n
MM13 cn c VDD VDD pch_mac W=0.2u L=30.00n
MM15 net20 cn net31 VDD pch_mac W=0.2u L=30.00n
MM19 net87 net16 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net31 c net87 VDD pch_mac W=120.00n L=30.00n
MM21 net16 net31 VDD VDD pch_mac W=200.00n L=30.00n
MM23 Q net16 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS NDQV4
.SUBCKT NDRNQV4 CKN D Q RDN VDD VSS
MM21 net164 net159 VDD VDD pch_mac W=200.00n L=30.00n
MM23 Q net164 VDD VDD pch_mac W=0.4u L=30.00n
MM11 c CKN VDD VDD pch_mac W=0.2u L=30.00n
MM1 net132 D VDD VDD pch_mac W=0.2u L=30.00n
MM19 net99 net164 VDD VDD pch_mac W=120.00n L=30.00n
MM8 net124 net144 VDD VDD pch_mac W=120.00n L=30.00n
MM26 net164 RDN VDD VDD pch_mac W=200.00n L=30.00n
MM0 net132 c net131 VDD pch_mac W=0.2u L=30.00n
MM15 net144 cn net159 VDD pch_mac W=0.2u L=30.00n
MM5 net144 net131 VDD VDD pch_mac W=200.00n L=30.00n
MM20 net159 c net99 VDD pch_mac W=120.00n L=30.00n
MM13 cn c VDD VDD pch_mac W=0.2u L=30.00n
MM7 net131 cn net124 VDD pch_mac W=0.2u L=30.00n
MM25 net124 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM3 net132 cn net131 VSS nch_mac W=0.12u L=30.00n
MM27 net168 net159 VSS VSS nch_mac W=0.2u L=30.00n
MM18 net164 RDN net168 VSS nch_mac W=0.2u L=30.00n
MM10 c CKN VSS VSS nch_mac W=0.2u L=30.00n
MM12 cn c VSS VSS nch_mac W=0.2u L=30.00n
MM17 net159 cn net152 VSS nch_mac W=120.00n L=30.00n
MM9 net176 net144 net180 VSS nch_mac W=120.00n L=30.00n
MM6 net131 c net176 VSS nch_mac W=120.00n L=30.00n
MM2 net132 D VSS VSS nch_mac W=0.2u L=30.00n
MM4 net144 net131 VSS VSS nch_mac W=0.2u L=30.00n
MM16 net152 net164 VSS VSS nch_mac W=120.00n L=30.00n
MM22 Q net164 VSS VSS nch_mac W=0.4u L=30.00n
MM24 net180 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM14 net144 c net159 VSS nch_mac W=0.2u L=30.00n
.ENDS NDRNQV4
.SUBCKT NDSRNQV4 CKN D Q RDN SDN VDD VSS
MM8 net165 cn net122 VDD pch_mac W=120.00n L=30.00n
MM24 net174 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM5 net174 net165 VDD VDD pch_mac W=200.00n L=30.00n
MM1 net170 D VDD VDD pch_mac W=120.00n L=30.00n
MM15 net174 cn net169 VDD pch_mac W=200.00n L=30.00n
MM0 net170 c net165 VDD pch_mac W=120.00n L=30.00n
MM20 net169 c net138 VDD pch_mac W=120.00n L=30.00n
MM37 net138 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM21 net198 net169 VDD VDD pch_mac W=200.00n L=30.00n
MM19 net138 net198 VDD VDD pch_mac W=120.00n L=30.00n
MM27 net198 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM13 cn c VDD VDD pch_mac W=200.00n L=30.00n
MM36 net122 net174 VDD VDD pch_mac W=120.00n L=30.00n
MM11 c CKN VDD VDD pch_mac W=200.00n L=30.00n
MM23 Q net198 VDD VDD pch_mac W=400.00n L=30.00n
MM35 net122 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM7 net165 c net194 VSS nch_mac W=120.00n L=30.00n
MM30 net202 net169 VSS VSS nch_mac W=200.00n L=30.00n
MM18 net198 RDN net202 VSS nch_mac W=200.00n L=30.00n
MM9 net194 net174 net186 VSS nch_mac W=120.00n L=30.00n
MM6 net186 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM26 net182 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM22 Q net198 VSS VSS nch_mac W=400.00n L=30.00n
MM4 net174 net165 net182 VSS nch_mac W=200.00n L=30.00n
MM14 net174 c net169 VSS nch_mac W=200.00n L=30.00n
MM3 net170 cn net165 VSS nch_mac W=120.00n L=30.00n
MM29 net158 SDN VSS VSS nch_mac W=120.00n L=30.00n
MM10 c CKN VSS VSS nch_mac W=200.00n L=30.00n
MM12 cn c VSS VSS nch_mac W=200.00n L=30.00n
MM2 net170 D VSS VSS nch_mac W=120.00n L=30.00n
MM16 net146 net198 net158 VSS nch_mac W=120.00n L=30.00n
MM17 net169 cn net146 VSS nch_mac W=120.00n L=30.00n
.ENDS NDSRNQV4
.SUBCKT NOR2V4 A1 A2 ZN VDD VSS
MMN1 ZN A1 VSS VSS nch_mac w=0.14u L=30.00n
MM0 ZN A2 VSS VSS nch_mac w=0.14u L=30.00n
MMP1 net15 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM1 ZN A1 net15 VDD pch_mac W=0.4u L=30.00n
.ENDS NOR2V4
.SUBCKT NOR2XBV4 A1 B1 ZN VDD VSS
MMN1 ZN net027 VSS VSS nch_mac W=0.4u L=30.00n
MM0 ZN B1 VSS VSS nch_mac W=0.4u L=30.00n
MM2 net027 A1 VSS VSS nch_mac W=0.19u L=30.00n
MMP1 net23 net027 VDD VDD pch_mac W=0.4u L=30.00n
MM3 net027 A1 VDD VDD pch_mac W=0.175u L=30.00n
MM1 ZN B1 net23 VDD pch_mac W=0.4u L=30.00n
.ENDS NOR2XBV4
.SUBCKT NOR3BBV4 A1 A2 B ZN VDD VSS
MM3 ZN A1N VSS VSS nch_mac W=0.38u L=30.00n
MM5 A1N A1 VSS VSS nch_mac W=0.175u L=30.00n
MM8 A2N A2 VSS VSS nch_mac W=0.175u L=30.00n
MM2 ZN B VSS VSS nch_mac W=0.4u L=30.00n
MM0 ZN A2N VSS VSS nch_mac W=0.38u L=30.00n
MM6 A2N A2 VDD VDD pch_mac W=0.175u L=30.00n
MM7 A1N A1 VDD VDD pch_mac W=0.175u L=30.00n
MM1 ZN A1N net24 VDD pch_mac W=0.4u L=30.00n
MM9 net051 B VDD VDD pch_mac W=0.4u L=30.00n
MM4 net24 A2N net051 VDD pch_mac W=0.4u L=30.00n
.ENDS NOR3BBV4
.SUBCKT NOR3V4 A1 A2 A3 ZN VDD VSS
MMN1 ZN A1 VSS VSS nch_mac W=0.24u L=30.00n
MM0 ZN A2 VSS VSS nch_mac W=0.24u L=30.00n
MM3 ZN A3 VSS VSS nch_mac W=0.24u L=30.00n
MMP1 net20 A2 net24 VDD pch_mac W=0.4u L=30.00n
MM1 ZN A1 net20 VDD pch_mac W=0.4u L=30.00n
MM2 net24 A3 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS NOR3V4
.SUBCKT NOR4BBV4 A1 A2 B1 B2 ZN VDD VSS
MM8 net89 A2 VSS VSS nch_mac W=200.00n L=30.00n
MM2 ZN B2 VSS VSS nch_mac W=400.00n L=30.00n
MM0 ZN B1 VSS VSS nch_mac W=400.00n L=30.00n
MM4 ZN net61 VSS VSS nch_mac W=400.00n L=30.00n
MM6 net61 A1 net89 VSS nch_mac W=200.00n L=30.00n
MM5 net61 A2 VDD VDD pch_mac W=200.00n L=30.00n
MM9 net72 B1 net60 VDD pch_mac W=400.00n L=30.00n
MM1 ZN net61 net72 VDD pch_mac W=400.00n L=30.00n
MM7 net61 A1 VDD VDD pch_mac W=200.00n L=30.00n
MM3 net60 B2 VDD VDD pch_mac W=400.00n L=30.00n
.ENDS NOR4BBV4
.SUBCKT NOR4V4 A1 A2 A3 A4 ZN VDD VSS
MMN1 ZN A1 VSS VSS nch_mac W=0.24u L=30.00n
MM0 ZN A2 VSS VSS nch_mac W=0.24u L=30.00n
MM3 ZN A3 VSS VSS nch_mac W=0.24u L=30.00n
MM4 ZN A4 VSS VSS nch_mac W=0.24u L=30.00n
MMP1 net25 A2 net29 VDD pch_mac W=0.39u L=30.00n
MM1 ZN A1 net25 VDD pch_mac W=0.39u L=30.00n
MM2 net29 A3 net33 VDD pch_mac W=0.39u L=30.00n
MM5 net33 A4 VDD VDD pch_mac W=0.39u L=30.00n
.ENDS NOR4V4
.SUBCKT NOR4XXBBV4 A1 A2 B1 B2 ZN VDD VSS
MM1 ZN B1 net38 VDD pch_mac W=0.4u L=30.00n
MM7 net27 A1 VDD VDD pch_mac W=0.175u L=30.00n
MM5 net27 A2 VDD VDD pch_mac W=0.175u L=30.00n
MM9 net38 B2 net26 VDD pch_mac W=0.4u L=30.00n
MM3 net26 net27 VDD VDD pch_mac W=0.4u L=30.00n
MM8 net55 A2 VSS VSS nch_mac W=0.175u L=30.00n
MM2 ZN B2 VSS VSS nch_mac W=0.4u L=30.00n
MM0 ZN B1 VSS VSS nch_mac W=0.4u L=30.00n
MM4 ZN net27 VSS VSS nch_mac W=0.4u L=30.00n
MM6 net27 A1 net55 VSS nch_mac W=0.175u L=30.00n
.ENDS NOR4XXBBV4
.SUBCKT OA112V4 A1 A2 B C Z VDD VSS
MM6 net30 B net14 VSS nch_mac W=0.2u L=30.00n
MM5 net14 C VSS VSS nch_mac W=0.2u L=30.00n
MM2 net043 A1 net30 VSS nch_mac W=0.2u L=30.00n
MM0 net043 A2 net30 VSS nch_mac W=0.2u L=30.00n
MM8 Z net043 VSS VSS nch_mac W=0.4u L=30.00n
MM4 net043 C VDD VDD pch_mac W=0.2u L=30.00n
MM3 net33 A2 VDD VDD pch_mac W=0.2u L=30.00n
MM9 net043 A1 net33 VDD pch_mac W=0.2u L=30.00n
MM7 Z net043 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net043 B VDD VDD pch_mac W=0.2u L=30.00n
.ENDS OA112V4
.SUBCKT OA12V4 A1 A2 B Z VDD VSS
MM0 Z net29 VSS VSS nch_mac W=0.4u L=30.00n
MM8 net027 B VSS VSS nch_mac W=0.2u L=30.00n
MM6 net29 A2 net027 VSS nch_mac W=0.2u L=30.00n
MM5 net29 A1 net027 VSS nch_mac W=0.2u L=30.00n
MM3 Z net29 VDD VDD pch_mac W=0.4u L=30.00n
MM7 net29 B VDD VDD pch_mac W=0.2u L=30.00n
MM4 net32 A2 VDD VDD pch_mac W=0.2u L=30.00n
MM1 net29 A1 net32 VDD pch_mac W=0.2u L=30.00n
.ENDS OA12V4
.SUBCKT OA13V4 A1 A2 A3 B Z VDD VSS
MM0 net26 A2 net30 VDD pch_mac W=0.2u L=30.00n
MM1 net51 B VDD VDD pch_mac W=0.2u L=30.00n
MM7 net51 A1 net26 VDD pch_mac W=0.2u L=30.00n
MM9 Z net51 VDD VDD pch_mac W=0.4u L=30.00n
MM3 net30 A3 VDD VDD pch_mac W=0.2u L=30.00n
MM5 net51 A1 net55 VSS nch_mac W=0.2u L=30.00n
MM8 net55 B VSS VSS nch_mac W=0.2u L=30.00n
MM2 net51 A3 net55 VSS nch_mac W=0.2u L=30.00n
MM4 Z net51 VSS VSS nch_mac W=0.4u L=30.00n
MM6 net51 A2 net55 VSS nch_mac W=0.2u L=30.00n
.ENDS OA13V4
.SUBCKT OA1B2V4 A1 A2 B Z VDD VSS
MMN1 Z net041 VSS VSS nch_mac W=0.4u L=30.00n
MM0 Z B VSS VSS nch_mac W=0.4u L=30.00n
MM2 net041 A2 VSS VSS nch_mac W=0.175u L=30.00n
MM3 net041 A1 VSS VSS nch_mac W=0.175u L=30.00n
MMP1 net28 net041 VDD VDD pch_mac W=0.4u L=30.00n
MM1 Z B net28 VDD pch_mac W=0.4u L=30.00n
MM5 net24 A2 VDD VDD pch_mac W=0.175u L=30.00n
MM4 net041 A1 net24 VDD pch_mac W=0.175u L=30.00n
.ENDS OA1B2V4
.SUBCKT OA212V4 A1 A2 B1 B2 C Z VDD VSS
MM11 Z net32 VSS VSS nch_mac W=400.00n L=30.00n
MM9 net55 C net64 VSS nch_mac W=0.2u L=30.00n
MM6 net64 B1 VSS VSS nch_mac W=0.2u L=30.00n
MM7 net64 B2 VSS VSS nch_mac W=0.2u L=30.00n
MM10 net32 A1 net55 VSS nch_mac W=0.2u L=30.00n
MM8 net32 A2 net55 VSS nch_mac W=0.2u L=30.00n
MM5 Z net32 VDD VDD pch_mac W=400.00n L=30.00n
MM0 net32 C VDD VDD pch_mac W=0.2u L=30.00n
MM4 net43 A2 VDD VDD pch_mac W=0.2u L=30.00n
MM3 net32 A1 net43 VDD pch_mac W=0.2u L=30.00n
MM2 net32 B1 net39 VDD pch_mac W=0.2u L=30.00n
MM1 net39 B2 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS OA212V4
.SUBCKT OA222V4 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM1 net48 B2 VDD VDD pch_mac W=0.19u L=30.00n
MM5 Z net41 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net41 C1 net44 VDD pch_mac W=0.19u L=30.00n
MM4 net52 A2 VDD VDD pch_mac W=0.19u L=30.00n
MM3 net41 A1 net52 VDD pch_mac W=0.19u L=30.00n
MM2 net41 B1 net48 VDD pch_mac W=0.19u L=30.00n
MM12 net44 C2 VDD VDD pch_mac W=0.19u L=30.00n
MM13 net41 A1 net69 VSS nch_mac W=0.175u L=30.00n
MM9 net41 A2 net69 VSS nch_mac W=0.175u L=30.00n
MM7 net69 B2 net77 VSS nch_mac W=0.175u L=30.00n
MM10 net77 C1 VSS VSS nch_mac W=0.175u L=30.00n
MM8 net77 C2 VSS VSS nch_mac W=0.175u L=30.00n
MM11 Z net41 VSS VSS nch_mac W=0.4u L=30.00n
MM6 net69 B1 net77 VSS nch_mac W=0.175u L=30.00n
.ENDS OA222V4
.SUBCKT OA22V4 A1 A2 B1 B2 Z VDD VSS
MM5 Z net42 VDD VDD pch_mac W=0.4u L=30.00n
MM4 net37 A2 VDD VDD pch_mac W=0.2u L=30.00n
MM1 net25 B2 VDD VDD pch_mac W=0.2u L=30.00n
MM3 net42 A1 net37 VDD pch_mac W=0.2u L=30.00n
MM2 net42 B1 net25 VDD pch_mac W=0.2u L=30.00n
MM11 Z net42 VSS VSS nch_mac W=0.4u L=30.00n
MM10 net54 B1 VSS VSS nch_mac W=0.2u L=30.00n
MM7 net42 A2 net54 VSS nch_mac W=0.2u L=30.00n
MM8 net54 B2 VSS VSS nch_mac W=0.2u L=30.00n
MM6 net42 A1 net54 VSS nch_mac W=0.2u L=30.00n
.ENDS OA22V4
.SUBCKT OA32V4 A1 A2 A3 B1 B2 Z VDD VSS
MM10 Z net27 VSS VSS nch_mac W=400.0n L=30.00n
MM9 net27 B2 net15 VSS nch_mac W=200.0n L=30.00n
MM2 net15 A3 VSS VSS nch_mac W=200.0n L=30.00n
MM5 net15 A1 VSS VSS nch_mac W=200.0n L=30.00n
MM6 net15 A2 VSS VSS nch_mac W=200.0n L=30.00n
MM8 net27 B1 net15 VSS nch_mac W=200.0n L=30.00n
MM11 Z net27 VDD VDD pch_mac W=400.0n L=30.00n
MM4 net38 B2 VDD VDD pch_mac W=200.0n L=30.00n
MM3 net50 A3 VDD VDD pch_mac W=200.0n L=30.00n
MM0 net42 A2 net50 VDD pch_mac W=200.0n L=30.00n
MM7 net27 A1 net42 VDD pch_mac W=200.0n L=30.00n
MM1 net27 B1 net38 VDD pch_mac W=200.0n L=30.00n
.ENDS OA32V4
.SUBCKT OA33V4 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM13 net36 A3 net52 VSS nch_mac W=0.2u L=30.00n
MM9 net36 A2 net52 VSS nch_mac W=0.2u L=30.00n
MM8 net36 A1 net52 VSS nch_mac W=0.2u L=30.00n
MM10 Z net36 VSS VSS nch_mac W=0.4u L=30.00n
MM2 net52 B3 VSS VSS nch_mac W=0.2u L=30.00n
MM6 net52 B2 VSS VSS nch_mac W=0.2u L=30.00n
MM5 net52 B1 VSS VSS nch_mac W=0.2u L=30.00n
MM12 net27 B3 VDD VDD pch_mac W=0.2u L=30.00n
MM3 net15 A3 VDD VDD pch_mac W=0.2u L=30.00n
MM0 net19 A2 net15 VDD pch_mac W=0.2u L=30.00n
MM4 net31 B2 net27 VDD pch_mac W=0.2u L=30.00n
MM7 net36 A1 net19 VDD pch_mac W=0.2u L=30.00n
MM1 net36 B1 net31 VDD pch_mac W=0.2u L=30.00n
MM11 Z net36 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS OA33V4
.SUBCKT OAI112V4 A1 A2 B C ZN VDD VSS
MM5 ZN C VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 net31 VDD pch_mac W=0.4u L=30.00n
MM4 ZN B VDD VDD pch_mac W=0.4u L=30.00n
MM0 net31 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM2 net43 B net52 VSS nch_mac W=0.4u L=30.00n
MM3 net52 C VSS VSS nch_mac W=0.4u L=30.00n
MMN1 ZN A2 net43 VSS nch_mac W=0.4u L=30.00n
MM1 ZN A1 net43 VSS nch_mac W=0.4u L=30.00n
.ENDS OAI112V4
.SUBCKT OAI12V4 A1 A2 B ZN VDD VSS
MM0 net32 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM4 ZN B VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 net32 VDD pch_mac W=0.4u L=30.00n
MM2 net36 B VSS VSS nch_mac W=0.4u L=30.00n
MMN1 ZN A1 net36 VSS nch_mac W=0.4u L=30.00n
MM1 ZN A2 net36 VSS nch_mac W=0.4u L=30.00n
.ENDS OAI12V4
.SUBCKT OAI13V4 A1 A2 A3 B ZN VDD VSS
MM0 net45 A2 net41 VDD pch_mac W=0.4u L=30.00n
MM8 net41 A3 VDD VDD pch_mac W=0.4u L=30.00n
MM4 ZN B VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 net45 VDD pch_mac W=0.4u L=30.00n
MMN1 ZN A2 net53 VSS nch_mac W=0.4u L=30.00n
MM1 ZN A3 net53 VSS nch_mac W=0.4u L=30.00n
MM2 net53 B VSS VSS nch_mac W=0.4u L=30.00n
MM9 ZN A1 net53 VSS nch_mac W=0.4u L=30.00n
.ENDS OAI13V4
.SUBCKT OAI212V4 A1 A2 B1 B2 C ZN VDD VSS
MM5 ZN C VDD VDD pch_mac W=0.4u L=30.00n
MM8 net41 B2 VDD VDD pch_mac W=0.4u L=30.00n
MMP1 ZN A1 net53 VDD pch_mac W=0.4u L=30.00n
MM0 net53 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM4 ZN B1 net41 VDD pch_mac W=0.4u L=30.00n
MMN1 net58 B2 VSS VSS nch_mac W=0.4u L=30.00n
MM1 net58 B1 VSS VSS nch_mac W=0.4u L=30.00n
MM3 net73 C net58 VSS nch_mac W=0.4u L=30.00n
MM9 ZN A2 net73 VSS nch_mac W=0.4u L=30.00n
MM2 ZN A1 net73 VSS nch_mac W=0.4u L=30.00n
.ENDS OAI212V4
.SUBCKT OAI21BV4 A B1 B2 ZN VDD VSS
MM5 net9 B1 VSS VSS nch_mac W=0.4u L=30.00n
MM6 net9 B2 VSS VSS nch_mac W=0.4u L=30.00n
MM8 ZN net17 net9 VSS nch_mac W=0.4u L=30.00n
MM0 net17 A VSS VSS nch_mac W=0.175u L=30.00n
MM1 ZN B1 net24 VDD pch_mac W=0.4u L=30.00n
MM4 net24 B2 VDD VDD pch_mac W=0.4u L=30.00n
MM7 ZN net17 VDD VDD pch_mac W=400.00n L=30.00n
MM3 net17 A VDD VDD pch_mac W=0.175u L=30.00n
.ENDS OAI21BV4
.SUBCKT OAI222V4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MMN1 ZN A2 net20 VSS nch_mac W=0.4u L=30.00n
MM1 ZN A1 net20 VSS nch_mac W=0.4u L=30.00n
MM3 net12 C1 VSS VSS nch_mac W=0.4u L=30.00n
MM2 net20 B1 net12 VSS nch_mac W=0.4u L=30.00n
MM9 net20 B2 net12 VSS nch_mac W=0.4u L=30.00n
MM12 net12 C2 VSS VSS nch_mac W=0.4u L=30.00n
MMP1 ZN A1 net43 VDD pch_mac W=0.4u L=30.00n
MM0 net43 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM4 ZN B1 net39 VDD pch_mac W=0.4u L=30.00n
MM11 ZN C1 net35 VDD pch_mac W=0.4u L=30.00n
MM10 net35 C2 VDD VDD pch_mac W=0.4u L=30.00n
MM8 net39 B2 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS OAI222V4
.SUBCKT OAI22BBV4 A1 A2 B1 B2 ZN VDD VSS
MMN1 net6 A2 VSS VSS nch_mac W=0.175u L=30.00n
MM1 net30 A1 net6 VSS nch_mac W=0.175u L=30.00n
MM3 ZN B1 net054 VSS nch_mac W=0.435u L=30.00n
MM2 net054 net30 VSS VSS nch_mac W=0.4u L=30.00n
MM6 ZN B2 net054 VSS nch_mac W=0.4u L=30.00n
MMP1 net30 A1 VDD VDD pch_mac W=0.175u L=30.00n
MM0 net30 A2 VDD VDD pch_mac W=0.175u L=30.00n
MM7 net37 B2 VDD VDD pch_mac W=0.4u L=30.00n
MM5 ZN net30 VDD VDD pch_mac W=0.4u L=30.00n
MM4 ZN B1 net37 VDD pch_mac W=0.435u L=30.00n
.ENDS OAI22BBV4
.SUBCKT OAI22V4 A1 A2 B1 B2 ZN VDD VSS
MMN1 ZN A2 net10 VSS nch_mac W=0.4u L=30.00n
MM1 ZN A1 net10 VSS nch_mac W=0.4u L=30.00n
MM2 net10 B1 VSS VSS nch_mac W=0.4u L=30.00n
MM9 net10 B2 VSS VSS nch_mac W=0.4u L=30.00n
MMP1 ZN A1 net29 VDD pch_mac W=0.4u L=30.00n
MM0 net29 A2 VDD VDD pch_mac W=0.4u L=30.00n
MM4 ZN B1 net25 VDD pch_mac W=0.4u L=30.00n
MM8 net25 B2 VDD VDD pch_mac W=0.4u L=30.00n
.ENDS OAI22V4
.SUBCKT OAI32V4 A1 A2 A3 B1 B2 ZN VDD VSS
MM8 ZN B1 net43 VSS nch_mac W=400.00n L=30.00n
MM6 net43 A2 VSS VSS nch_mac W=400.00n L=30.00n
MM5 net43 A1 VSS VSS nch_mac W=400.00n L=30.00n
MM2 net43 A3 VSS VSS nch_mac W=400.00n L=30.00n
MM9 ZN B2 net43 VSS nch_mac W=400.00n L=30.00n
MM1 ZN B1 net10 VDD pch_mac W=400.00n L=30.00n
MM7 ZN A1 net14 VDD pch_mac W=400.00n L=30.00n
MM0 net14 A2 net18 VDD pch_mac W=400.00n L=30.00n
MM3 net18 A3 VDD VDD pch_mac W=400.00n L=30.00n
MM4 net10 B2 VDD VDD pch_mac W=400.00n L=30.00n
.ENDS OAI32V4
.SUBCKT OAI33V4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM11 net041 A2 VSS VSS nch_mac W=400.00n L=30.00n
MM2 net041 A1 VSS VSS nch_mac W=400.00n L=30.00n
MM9 ZN B3 net041 VSS nch_mac W=400.00n L=30.00n
MM1 ZN B1 net041 VSS nch_mac W=400.00n L=30.00n
MM13 net041 A3 VSS VSS nch_mac W=400.00n L=30.00n
MMN1 ZN B2 net041 VSS nch_mac W=400.00n L=30.00n
MM12 net076 B3 VDD VDD pch_mac W=400.00n L=30.00n
MM4 ZN B1 net071 VDD pch_mac W=400.00n L=30.00n
MM8 net065 A3 VDD VDD pch_mac W=400.00n L=30.00n
MM10 net071 B2 net076 VDD pch_mac W=400.00n L=30.00n
MM0 net067 A2 net065 VDD pch_mac W=400.00n L=30.00n
MMP1 ZN A1 net067 VDD pch_mac W=400.00n L=30.00n
.ENDS OAI33V4
.SUBCKT OR2V4 A1 A2 Z VDD VSS
MMN1 net12 A1 VSS VSS nch_mac W=0.2u L=30.00n
MM2 Z net12 VSS VSS nch_mac W=0.4u L=30.00n
MM0 net12 A2 VSS VSS nch_mac W=0.2u L=30.00n
MMP1 net23 A2 VDD VDD pch_mac W=0.2u L=30.00n
MM4 Z net12 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net12 A1 net23 VDD pch_mac W=0.2u L=30.00n
.ENDS OR2V4
.SUBCKT OR3V4 A1 A2 A3 Z VDD VSS
MMP1 net20 A2 net8 VDD pch_mac W=0.2u L=30.00n
MM5 net8 A3 VDD VDD pch_mac W=0.2u L=30.00n
MM4 Z net21 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net21 A1 net20 VDD pch_mac W=0.2u L=30.00n
MMN1 net21 A1 VSS VSS nch_mac W=0.2u L=30.00n
MM2 Z net21 VSS VSS nch_mac W=0.4u L=30.00n
MM0 net21 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM3 net21 A3 VSS VSS nch_mac W=0.2u L=30.00n
.ENDS OR3V4
.SUBCKT OR4V4 A1 A2 A3 A4 Z VDD VSS
MM7 net6 A1 VSS VSS nch_mac W=0.2u L=30.00n
MM3 net6 A4 VSS VSS nch_mac W=0.2u L=30.00n
MM0 net6 A3 VSS VSS nch_mac W=0.2u L=30.00n
MM2 Z net6 VSS VSS nch_mac W=0.4u L=30.00n
MMN1 net6 A2 VSS VSS nch_mac W=0.2u L=30.00n
MM1 net6 A1 net33 VDD pch_mac W=0.2u L=30.00n
MM4 Z net6 VDD VDD pch_mac W=0.4u L=30.00n
MM5 net45 A3 net41 VDD pch_mac W=0.2u L=30.00n
MMP1 net33 A2 net45 VDD pch_mac W=0.2u L=30.00n
MM6 net41 A4 VDD VDD pch_mac W=0.2u L=30.00n
.ENDS OR4V4
.SUBCKT SDGRNQNV4 CK D QN RN SE SI VDD VSS
MM18 net129 net96 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net96 cn net113 VSS nch_mac W=120.00n L=30.00n
MM9 net121 net137 VSS VSS nch_mac W=120.00n L=30.00n
MM3 net149 cn net120 VSS nch_mac W=200.00n L=30.00n
MM16 net113 net129 VSS VSS nch_mac W=120.00n L=30.00n
MM31 net149 SE net141 VSS nch_mac W=120.00n L=30.00n
MM22 QN net96 VSS VSS nch_mac W=400.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=120.00n L=30.00n
MM14 net137 c net96 VSS nch_mac W=200.00n L=30.00n
MM34 net149 D net81 VSS nch_mac W=200.00n L=30.00n
MM32 net85 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM33 net81 RN net85 VSS nch_mac W=200.00n L=30.00n
MM6 net120 c net121 VSS nch_mac W=120.00n L=30.00n
MM30 net141 SI VSS VSS nch_mac W=120.00n L=30.00n
MM4 net137 net120 VSS VSS nch_mac W=200.00n L=30.00n
MM25 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM23 QN net96 VDD VDD pch_mac W=400.00n L=30.00n
MM20 net96 c net192 VDD pch_mac W=120.00n L=30.00n
MM21 net129 net96 VDD VDD pch_mac W=120.00n L=30.00n
MM0 net149 c net120 VDD pch_mac W=200.00n L=30.00n
MM28 net164 SI VDD VDD pch_mac W=120.00n L=30.00n
MM8 net216 net137 VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=120.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=120.00n L=30.00n
MM5 net137 net120 VDD VDD pch_mac W=200.00n L=30.00n
MM19 net192 net129 VDD VDD pch_mac W=120.00n L=30.00n
MM15 net137 cn net96 VDD pch_mac W=200.00n L=30.00n
MM24 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM29 net149 SEN net164 VDD pch_mac W=120.00n L=30.00n
MM37 net152 SE VDD VDD pch_mac W=200.00n L=30.00n
MM36 net149 RN net152 VDD pch_mac W=200.00n L=30.00n
MM7 net120 cn net216 VDD pch_mac W=120.00n L=30.00n
MM35 net149 D net152 VDD pch_mac W=200.00n L=30.00n
.ENDS SDGRNQNV4
.SUBCKT SDGRSNQNV4 CK D QN RN SE SI SN VDD VSS
MM9 net139 net155 VSS VSS nch_mac W=120.00n L=30.00n
MM3 net103 cn net138 VSS nch_mac W=200.00n L=30.00n
MM16 net131 net147 VSS VSS nch_mac W=120.00n L=30.00n
MM31 net103 SE net159 VSS nch_mac W=120.00n L=30.00n
MM22 QN net114 VSS VSS nch_mac W=400.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM14 net155 c net114 VSS nch_mac W=200.00n L=30.00n
MM38 net103 snn net95 VSS nch_mac W=120.00n L=30.00n
MM2 net103 D net95 VSS nch_mac W=200.00n L=30.00n
MM26 net99 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM33 net95 RN net99 VSS nch_mac W=200.00n L=30.00n
MM35 snn SN VSS VSS nch_mac W=120.00n L=30.00n
MM6 net138 c net139 VSS nch_mac W=120.00n L=30.00n
MM30 net159 SI VSS VSS nch_mac W=120.00n L=30.00n
MM4 net155 net138 VSS VSS nch_mac W=200.00n L=30.00n
MM25 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM18 net147 net114 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net114 cn net131 VSS nch_mac W=120.00n L=30.00n
MM24 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM29 net103 SEN net190 VDD pch_mac W=120.00n L=30.00n
MM1 net103 D net186 VDD pch_mac W=200.00n L=30.00n
MM34 net103 RN net170 VDD pch_mac W=120.00n L=30.00n
MM36 snn SN VDD VDD pch_mac W=120.00n L=30.00n
MM27 net170 SE VDD VDD pch_mac W=200.00n L=30.00n
MM37 net186 snn net170 VDD pch_mac W=200.00n L=30.00n
MM7 net138 cn net242 VDD pch_mac W=120.00n L=30.00n
MM5 net155 net138 VDD VDD pch_mac W=200.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM19 net218 net147 VDD VDD pch_mac W=120.00n L=30.00n
MM0 net103 c net138 VDD pch_mac W=200.00n L=30.00n
MM23 QN net114 VDD VDD pch_mac W=400.00n L=30.00n
MM20 net114 c net218 VDD pch_mac W=120.00n L=30.00n
MM21 net147 net114 VDD VDD pch_mac W=120.00n L=30.00n
MM28 net190 SI VDD VDD pch_mac W=120.00n L=30.00n
MM8 net242 net155 VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM15 net155 cn net114 VDD pch_mac W=200.00n L=30.00n
.ENDS SDGRSNQNV4
.SUBCKT SDQNV4 CK D QN SE SI VDD VSS
MM1 net131 D net134 VDD pch_mac W=200.00n L=30.00n
MM27 net134 SE VDD VDD pch_mac W=200.00n L=30.00n
MM29 net131 SEN net126 VDD pch_mac W=0.2u L=30.00n
MM28 net126 SI VDD VDD pch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM23 QN net162 VDD VDD pch_mac W=0.4u L=30.00n
MM21 net167 net162 VDD VDD pch_mac W=120.00n L=30.00n
MM5 net163 net199 VDD VDD pch_mac W=0.2u L=30.00n
MM15 net163 cn net162 VDD pch_mac W=0.2u L=30.00n
MM20 net162 c net94 VDD pch_mac W=0.2u L=30.00n
MM7 net199 cn net90 VDD pch_mac W=120.00n L=30.00n
MM19 net94 net167 VDD VDD pch_mac W=0.2u L=30.00n
MM8 net90 net163 VDD VDD pch_mac W=120.00n L=30.00n
MM24 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM33 net199 c net131 VDD pch_mac W=0.2u L=30.00n
MM31 net191 SI net187 VSS nch_mac W=0.2u L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM25 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM32 net199 cn net191 VSS nch_mac W=0.2u L=30.00n
MM26 net195 D VSS VSS nch_mac W=200.00n L=30.00n
MM2 net191 SEN net195 VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM22 QN net162 VSS VSS nch_mac W=0.4u L=30.00n
MM18 net167 net162 VSS VSS nch_mac W=120.00n L=30.00n
MM4 net163 net199 VSS VSS nch_mac W=0.2u L=30.00n
MM30 net187 SE VSS VSS nch_mac W=0.2u L=30.00n
MM14 net163 c net162 VSS nch_mac W=0.2u L=30.00n
MM16 net155 net167 VSS VSS nch_mac W=0.2u L=30.00n
MM9 net151 net163 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net162 cn net155 VSS nch_mac W=0.2u L=30.00n
MM6 net199 c net151 VSS nch_mac W=120.00n L=30.00n
.ENDS SDQNV4
.SUBCKT SDQV4 CK D Q SE SI VDD VSS
MM32 net78 cn net86 VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM31 net86 SI net90 VSS nch_mac W=0.2u L=30.00n
MM26 net82 D VSS VSS nch_mac W=200.00n L=30.00n
MM2 net86 SEN net82 VSS nch_mac W=200.00n L=30.00n
MM22 Q net106 VSS VSS nch_mac W=0.4u L=30.00n
MM30 net90 SE VSS VSS nch_mac W=0.2u L=30.00n
MM4 net110 net78 VSS VSS nch_mac W=0.2u L=30.00n
MM25 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM6 net78 c net122 VSS nch_mac W=120.00n L=30.00n
MM17 net117 cn net118 VSS nch_mac W=120.00n L=30.00n
MM18 net106 net117 VSS VSS nch_mac W=0.2u L=30.00n
MM16 net118 net106 VSS VSS nch_mac W=120.00n L=30.00n
MM9 net122 net110 VSS VSS nch_mac W=120.00n L=30.00n
MM14 net110 c net117 VSS nch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM28 net157 SI VDD VDD pch_mac W=0.2u L=30.00n
MM7 net78 cn net189 VDD pch_mac W=120.00n L=30.00n
MM20 net117 c net185 VDD pch_mac W=120.00n L=30.00n
MM19 net185 net106 VDD VDD pch_mac W=120.00n L=30.00n
MM27 net149 SE VDD VDD pch_mac W=200.00n L=30.00n
MM21 net106 net117 VDD VDD pch_mac W=0.2u L=30.00n
MM33 net78 c net146 VDD pch_mac W=0.2u L=30.00n
MM5 net110 net78 VDD VDD pch_mac W=0.2u L=30.00n
MM29 net146 SEN net157 VDD pch_mac W=0.2u L=30.00n
MM8 net189 net110 VDD VDD pch_mac W=120.00n L=30.00n
MM23 Q net106 VDD VDD pch_mac W=0.4u L=30.00n
MM1 net146 D net149 VDD pch_mac W=200.00n L=30.00n
MM24 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM15 net110 cn net117 VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
.ENDS SDQV4
.SUBCKT SDRNQNV4 CK D QN RDN SE SI VDD VSS
MM3 QN net213 VDD VDD pch_mac W=400.00n L=30.00n
MM26 net189 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM15 net149 cn net200 VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM20 net213 c net200 VDD pch_mac W=120.00n L=30.00n
MM19 net213 net189 VDD VDD pch_mac W=200.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM34 SEN SE VDD VDD pch_mac W=120.0n L=30.00n
MM8 net125 net149 VDD VDD pch_mac W=120.00n L=30.00n
MM33 net177 c net93 VDD pch_mac W=0.2u L=30.00n
MM1 net93 D net96 VDD pch_mac W=200.00n L=30.00n
MM29 net96 SE VDD VDD pch_mac W=200.00n L=30.00n
MM5 net149 net177 VDD VDD pch_mac W=0.2u L=30.00n
MM36 net93 SEN net88 VDD pch_mac W=120.0n L=30.00n
MM21 net189 net200 VDD VDD pch_mac W=200.00n L=30.00n
MM37 net88 SI VDD VDD pch_mac W=120.0n L=30.00n
MM7 net177 cn net125 VDD pch_mac W=0.2u L=30.00n
MM25 net125 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM31 net201 SI net161 VSS nch_mac W=120.0n L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM30 net161 SE VSS VSS nch_mac W=120.0n L=30.00n
MM9 net157 net149 net173 VSS nch_mac W=120.00n L=30.00n
MM6 net177 c net157 VSS nch_mac W=120.00n L=30.00n
MM24 net173 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM32 net177 cn net201 VSS nch_mac W=200.00n L=30.00n
MM4 net149 net177 VSS VSS nch_mac W=0.2u L=30.00n
MM27 net205 net200 VSS VSS nch_mac W=200.00n L=30.00n
MM35 SEN SE VSS VSS nch_mac W=120.0n L=30.00n
MM17 net213 cn net200 VSS nch_mac W=120.00n L=30.00n
MM0 QN net213 VSS VSS nch_mac W=400.00n L=30.00n
MM16 net213 net189 VSS VSS nch_mac W=200.00n L=30.00n
MM2 net201 SEN net181 VSS nch_mac W=200.00n L=30.00n
MM14 net149 c net200 VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM18 net189 RDN net205 VSS nch_mac W=200.00n L=30.00n
MM28 net181 D VSS VSS nch_mac W=200.00n L=30.00n
.ENDS SDRNQNV4
.SUBCKT SDRNQV4 CK D Q RDN SE SI VDD VSS
MM27 net119 net118 VSS VSS nch_mac W=0.2u L=30.00n
MM30 net87 SE VSS VSS nch_mac W=0.2u L=30.00n
MM22 Q net123 VSS VSS nch_mac W=0.4u L=30.00n
MM32 net99 cn net91 VSS nch_mac W=120.00n L=30.00n
MM17 net118 cn net135 VSS nch_mac W=120.00n L=30.00n
MM18 net123 RDN net119 VSS nch_mac W=0.2u L=30.00n
MM31 net91 SI net87 VSS nch_mac W=0.2u L=30.00n
MM2 net91 SEN net95 VSS nch_mac W=200.00n L=30.00n
MM14 net131 c net118 VSS nch_mac W=0.2u L=30.00n
MM28 net95 D VSS VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM35 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM16 net135 net123 VSS VSS nch_mac W=120.00n L=30.00n
MM4 net131 net99 VSS VSS nch_mac W=0.2u L=30.00n
MM9 net143 net131 net127 VSS nch_mac W=120.00n L=30.00n
MM6 net99 c net143 VSS nch_mac W=120.00n L=30.00n
MM24 net127 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM26 net123 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM25 net199 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM20 net118 c net214 VDD pch_mac W=120.00n L=30.00n
MM5 net131 net99 VDD VDD pch_mac W=0.2u L=30.00n
MM8 net199 net131 VDD VDD pch_mac W=120.00n L=30.00n
MM15 net131 cn net118 VDD pch_mac W=0.2u L=30.00n
MM34 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM21 net123 net118 VDD VDD pch_mac W=0.2u L=30.00n
MM29 net170 SE VDD VDD pch_mac W=200.00n L=30.00n
MM1 net167 D net170 VDD pch_mac W=200.00n L=30.00n
MM23 Q net123 VDD VDD pch_mac W=0.4u L=30.00n
MM19 net214 net123 VDD VDD pch_mac W=120.00n L=30.00n
MM37 net162 SI VDD VDD pch_mac W=0.2u L=30.00n
MM33 net99 c net167 VDD pch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=0.2u L=30.00n
MM7 net99 cn net199 VDD pch_mac W=0.2u L=30.00n
MM36 net167 SEN net162 VDD pch_mac W=0.2u L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
.ENDS SDRNQV4
.SUBCKT SDRQNV4 CK D QN RD SE SI VDD VSS
MM2 net139 D net119 VSS nch_mac W=200.00n L=30.00n
MM27 net146 RD VSS VSS nch_mac W=120.00n L=30.00n
MM31 net139 SE net107 VSS nch_mac W=120.00n L=30.00n
MM17 net146 cn net151 VSS nch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM0 net119 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM35 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM30 net107 SI VSS VSS nch_mac W=120.00n L=30.00n
MM6 net90 c net99 VSS nch_mac W=120.00n L=30.00n
MM9 net99 net91 VSS VSS nch_mac W=120.00n L=30.00n
MM22 QN net146 VSS VSS nch_mac W=400.00n L=30.00n
MM4 net91 net90 VSS VSS nch_mac W=200.00n L=30.00n
MM32 net139 cn net90 VSS nch_mac W=200.00n L=30.00n
MM18 net153 net146 VSS VSS nch_mac W=120.00n L=30.00n
MM16 net151 net153 VSS VSS nch_mac W=120.00n L=30.00n
MM25 net91 RD VSS VSS nch_mac W=120.00n L=30.00n
MM14 net91 c net146 VSS nch_mac W=200.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM28 net182 SI VDD VDD pch_mac W=120.00n L=30.00n
MM7 net90 cn net202 VDD pch_mac W=120.00n L=30.00n
MM8 net202 net91 VDD VDD pch_mac W=120.00n L=30.00n
MM19 net166 net153 net194 VDD pch_mac W=120.00n L=30.00n
MM3 net174 SE VDD VDD pch_mac W=200.00n L=30.00n
MM21 net153 net146 VDD VDD pch_mac W=120.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM34 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM24 net162 RD VDD VDD pch_mac W=200.00n L=30.00n
MM33 net139 c net90 VDD pch_mac W=200.00n L=30.00n
MM29 net139 SEN net182 VDD pch_mac W=120.00n L=30.00n
MM26 net194 RD VDD VDD pch_mac W=120.00n L=30.00n
MM1 net139 D net174 VDD pch_mac W=200.00n L=30.00n
MM15 net91 cn net146 VDD pch_mac W=200.00n L=30.00n
MM20 net146 c net166 VDD pch_mac W=120.00n L=30.00n
MM5 net91 net90 net162 VDD pch_mac W=200.00n L=30.00n
MM23 QN net146 VDD VDD pch_mac W=400.00n L=30.00n
.ENDS SDRQNV4
.SUBCKT SDRQV4 CK D Q RD SE SI VDD VSS
MM18 net223 net0146 VSS VSS nch_mac W=200.00n L=30.00n
MM32 net233 cn net228 VSS nch_mac W=200.00n L=30.00n
MM4 net241 net228 VSS VSS nch_mac W=200.00n L=30.00n
MM22 Q net223 VSS VSS nch_mac W=400.00n L=30.00n
MM9 net213 net241 VSS VSS nch_mac W=120.00n L=30.00n
MM6 net228 c net213 VSS nch_mac W=120.00n L=30.00n
MM30 net265 SI VSS VSS nch_mac W=120.00n L=30.00n
MM35 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM0 net261 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM17 net0146 cn net221 VSS nch_mac W=120.00n L=30.00n
MM31 net233 SE net265 VSS nch_mac W=120.00n L=30.00n
MM27 net0146 RD VSS VSS nch_mac W=200.00n L=30.00n
MM2 net233 D net261 VSS nch_mac W=200.00n L=30.00n
MM14 net241 c net0146 VSS nch_mac W=200.00n L=30.00n
MM25 net241 RD VSS VSS nch_mac W=120.00n L=30.00n
MM16 net221 net223 VSS VSS nch_mac W=120.00n L=30.00n
MM23 Q net223 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net241 net228 net184 VDD pch_mac W=200.00n L=30.00n
MM20 net0146 c net152 VDD pch_mac W=120.00n L=30.00n
MM15 net241 cn net0146 VDD pch_mac W=200.00n L=30.00n
MM1 net233 D net176 VDD pch_mac W=200.00n L=30.00n
MM26 net148 RD VDD VDD pch_mac W=120.00n L=30.00n
MM29 net233 SEN net180 VDD pch_mac W=120.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM21 net223 net0146 VDD VDD pch_mac W=200.00n L=30.00n
MM19 net152 net223 net148 VDD pch_mac W=120.00n L=30.00n
MM8 net144 net241 VDD VDD pch_mac W=120.00n L=30.00n
MM7 net228 cn net144 VDD pch_mac W=120.00n L=30.00n
MM28 net180 SI VDD VDD pch_mac W=120.00n L=30.00n
MM33 net233 c net228 VDD pch_mac W=200.00n L=30.00n
MM34 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM24 net184 RD VDD VDD pch_mac W=200.00n L=30.00n
MM3 net176 SE VDD VDD pch_mac W=200.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
.ENDS SDRQV4
.SUBCKT SDSRNQV4 CK D Q RDN SDN SE SI VDD VSS
MM3 net148 cn net159 VSS nch_mac W=200.00n L=30.00n
MM14 net140 c net155 VSS nch_mac W=200.00n L=30.00n
MM34 net148 D net132 VSS nch_mac W=200.00n L=30.00n
MM1 net148 SE net128 VSS nch_mac W=120.00n L=30.00n
MM4 net140 net159 net120 VSS nch_mac W=200.00n L=30.00n
MM22 Q net100 VSS VSS nch_mac W=400.00n L=30.00n
MM33 net132 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM2 net128 SI VSS VSS nch_mac W=120.00n L=30.00n
MM44 net124 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM26 net120 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM43 net116 net140 net124 VSS nch_mac W=120.00n L=30.00n
MM9 net159 c net116 VSS nch_mac W=120.00n L=30.00n
MM39 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM30 net104 net155 VSS VSS nch_mac W=200.00n L=30.00n
MM18 net100 RDN net104 VSS nch_mac W=200.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=200.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=200.00n L=30.00n
MM17 net155 cn net164 VSS nch_mac W=120.00n L=30.00n
MM16 net164 net100 net160 VSS nch_mac W=120.00n L=30.00n
MM29 net160 SDN VSS VSS nch_mac W=120.00n L=30.00n
MM7 net232 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM27 net100 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM21 net100 net155 VDD VDD pch_mac W=200.00n L=30.00n
MM0 net148 c net159 VDD pch_mac W=200.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=200.00n L=30.00n
MM38 net148 D net215 VDD pch_mac W=200.00n L=30.00n
MM40 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM35 net148 SEN net211 VDD pch_mac W=120.00n L=30.00n
MM5 net140 net159 VDD VDD pch_mac W=200.00n L=30.00n
MM15 net140 cn net155 VDD pch_mac W=200.00n L=30.00n
MM23 Q net100 VDD VDD pch_mac W=400.00n L=30.00n
MM24 net140 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM36 net211 SI VDD VDD pch_mac W=120.00n L=30.00n
MM25 net180 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM19 net180 net100 VDD VDD pch_mac W=120.00n L=30.00n
MM6 net232 net140 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net155 c net180 VDD pch_mac W=120.00n L=30.00n
MM8 net159 cn net232 VDD pch_mac W=120.00n L=30.00n
MM37 net215 SE VDD VDD pch_mac W=200.00n L=30.00n
.ENDS SDSRNQV4
.SUBCKT SDSNQNV4 CK D QN SDN SE SI VDD VSS
MM28 net318 SDN VDD VDD pch_mac W=0.2u L=30.00n
MM7 net358 cn net241 VDD pch_mac W=120.00n L=30.00n
MM23 QN net345 VDD VDD pch_mac W=0.4u L=30.00n
MM33 net358 c net290 VDD pch_mac W=0.2u L=30.00n
MM1 net290 D net293 VDD pch_mac W=200.00n L=30.00n
MM29 net270 SDN VDD VDD pch_mac W=0.2u L=30.00n
MM20 net345 c net270 VDD pch_mac W=0.2u L=30.00n
MM5 net318 net358 VDD VDD pch_mac W=0.2u L=30.00n
MM19 net270 net324 VDD VDD pch_mac W=0.2u L=30.00n
MM36 net290 SEN net301 VDD pch_mac W=0.2u L=30.00n
MM0 net293 SE VDD VDD pch_mac W=200.00n L=30.00n
MM8 net241 net318 VDD VDD pch_mac W=120.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
MM21 net324 net345 VDD VDD pch_mac W=120.00n L=30.00n
MM15 net318 cn net345 VDD pch_mac W=0.2u L=30.00n
MM34 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM37 net301 SI VDD VDD pch_mac W=0.2u L=30.00n
MM3 net366 SEN net362 VSS nch_mac W=200.00n L=30.00n
MM9 net306 net318 VSS VSS nch_mac W=120.00n L=30.00n
MM2 net362 D VSS VSS nch_mac W=200.00n L=30.00n
MM6 net358 c net306 VSS nch_mac W=120.00n L=30.00n
MM17 net345 cn net330 VSS nch_mac W=0.2u L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM18 net324 net345 VSS VSS nch_mac W=120.00n L=30.00n
MM31 net366 SI net370 VSS nch_mac W=0.2u L=30.00n
MM30 net370 SE VSS VSS nch_mac W=0.2u L=30.00n
MM25 net322 net324 VSS VSS nch_mac W=0.2u L=30.00n
MM22 QN net345 VSS VSS nch_mac W=0.4u L=30.00n
MM24 net314 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM4 net318 net358 net314 VSS nch_mac W=200.00n L=30.00n
MM35 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM16 net330 SDN net322 VSS nch_mac W=0.2u L=30.00n
MM32 net358 cn net366 VSS nch_mac W=0.2u L=30.00n
MM14 net318 c net345 VSS nch_mac W=0.2u L=30.00n
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
.ENDS SDSNQNV4
.SUBCKT SDSNQV4 CK D Q SDN SE SI VDD VSS
MM10 cn CK VSS VSS nch_mac W=0.2u L=30.00n
MM30 net140 SE VSS VSS nch_mac W=0.2u L=30.00n
MM32 net76 cn net132 VSS nch_mac W=0.2u L=30.00n
MM12 c cn VSS VSS nch_mac W=0.2u L=30.00n
MM3 net132 SEN net104 VSS nch_mac W=200.00n L=30.00n
MM6 net76 c net124 VSS nch_mac W=120.00n L=30.00n
MM9 net124 net96 VSS VSS nch_mac W=120.00n L=30.00n
MM17 net83 cn net88 VSS nch_mac W=120.00n L=30.00n
MM31 net132 SI net140 VSS nch_mac W=0.2u L=30.00n
MM18 net90 net83 VSS VSS nch_mac W=0.2u L=30.00n
MM25 net108 SDN VSS VSS nch_mac W=120.00n L=30.00n
MM2 net104 D VSS VSS nch_mac W=200.00n L=30.00n
MM24 net100 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM4 net96 net76 net100 VSS nch_mac W=200.00n L=30.00n
MM22 Q net90 VSS VSS nch_mac W=0.4u L=30.00n
MM16 net88 net90 net108 VSS nch_mac W=120.00n L=30.00n
MM35 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM14 net96 c net83 VSS nch_mac W=0.2u L=30.00n
MM33 net76 c net212 VDD pch_mac W=0.2u L=30.00n
MM1 net212 D net215 VDD pch_mac W=200.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=0.2u L=30.00n
MM8 net199 net96 VDD VDD pch_mac W=120.00n L=30.00n
MM36 net212 SEN net207 VDD pch_mac W=0.2u L=30.00n
MM37 net207 SI VDD VDD pch_mac W=0.2u L=30.00n
MM7 net76 cn net199 VDD pch_mac W=120.00n L=30.00n
MM28 net96 SDN VDD VDD pch_mac W=0.2u L=30.00n
MM5 net96 net76 VDD VDD pch_mac W=0.2u L=30.00n
MM20 net83 c net160 VDD pch_mac W=120.00n L=30.00n
MM19 net160 net90 VDD VDD pch_mac W=120.00n L=30.00n
MM23 Q net90 VDD VDD pch_mac W=0.4u L=30.00n
MM0 net215 SE VDD VDD pch_mac W=200.00n L=30.00n
MM21 net90 net83 VDD VDD pch_mac W=0.2u L=30.00n
MM15 net96 cn net83 VDD pch_mac W=0.2u L=30.00n
MM29 net160 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM34 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
.ENDS SDSNQV4
.SUBCKT SEDRNQNV4 CK D E QN RDN SE SI VDD VSS
MM17 s cn net143 VSS nch_mac W=120.00n L=30.00n
MM31 net115 SE net187 VSS nch_mac W=120.00n L=30.00n
MM27 s R VSS VSS nch_mac W=120.00n L=30.00n
MM40 net155 s net122 VSS nch_mac W=120.00n L=30.00n
MM1 net115 en net155 VSS nch_mac W=120.00n L=30.00n
MM25 net131 R VSS VSS nch_mac W=120.00n L=30.00n
MM16 net143 net145 VSS VSS nch_mac W=120.00n L=30.00n
MM22 QN s VSS VSS nch_mac W=400.00n L=30.00n
MM14 net131 c s VSS nch_mac W=200.00n L=30.00n
MM4 net131 net130 VSS VSS nch_mac W=200.00n L=30.00n
MM32 net115 cn net130 VSS nch_mac W=200.00n L=30.00n
MM41 net122 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM39 net119 E net122 VSS nch_mac W=200.00n L=30.00n
MM38 net115 D net119 VSS nch_mac W=200.00n L=30.00n
MM18 net145 s VSS VSS nch_mac W=120.00n L=30.00n
MM36 R RDN VSS VSS nch_mac W=120.00n L=30.00n
MM9 net195 net131 VSS VSS nch_mac W=120.00n L=30.00n
MM6 net130 c net195 VSS nch_mac W=120.00n L=30.00n
MM30 net187 SI VSS VSS nch_mac W=120.00n L=30.00n
MM35 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM12 c cn VSS VSS nch_mac W=120.00n L=30.00n
MM0 en E VSS VSS nch_mac W=120.00n L=30.00n
MM10 cn CK VSS VSS nch_mac W=120.00n L=30.00n
MM34 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM2 net258 SE VDD VDD pch_mac W=200.00n L=30.00n
MM11 cn CK VDD VDD pch_mac W=120.00n L=30.00n
MM42 net115 D net262 VDD pch_mac W=200.00n L=30.00n
MM37 R RDN VDD VDD pch_mac W=120.00n L=30.00n
MM3 net262 en net258 VDD pch_mac W=200.00n L=30.00n
MM21 net145 s VDD VDD pch_mac W=120.00n L=30.00n
MM19 net290 net145 net238 VDD pch_mac W=120.00n L=30.00n
MM7 net130 cn net230 VDD pch_mac W=120.00n L=30.00n
MM8 net230 net131 VDD VDD pch_mac W=120.00n L=30.00n
MM28 net278 SI VDD VDD pch_mac W=120.00n L=30.00n
MM33 net115 c net130 VDD pch_mac W=200.00n L=30.00n
MM23 QN s VDD VDD pch_mac W=400.00n L=30.00n
MM5 net131 net130 net294 VDD pch_mac W=200.00n L=30.00n
MM15 net131 cn s VDD pch_mac W=200.00n L=30.00n
MM26 net238 R VDD VDD pch_mac W=120.00n L=30.00n
MM29 net115 SEN net278 VDD pch_mac W=120.00n L=30.00n
MM45 en E VDD VDD pch_mac W=120.00n L=30.00n
MM44 net115 E net270 VDD pch_mac W=120.00n L=30.00n
MM43 net270 s net258 VDD pch_mac W=120.00n L=30.00n
MM24 net294 R VDD VDD pch_mac W=200.00n L=30.00n
MM20 s c net290 VDD pch_mac W=120.00n L=30.00n
MM13 c cn VDD VDD pch_mac W=200.00n L=30.00n
.ENDS SEDRNQNV4
.SUBCKT SNDQV4 CKN D Q SE SI VDD VSS
MM11 c CKN VDD VDD pch_mac W=200.00n L=30.00n
MM0 net129 SE VDD VDD pch_mac W=200.00n L=30.00n
MM23 Q net146 VDD VDD pch_mac W=0.4u L=30.00n
MM13 cn c VDD VDD pch_mac W=0.2u L=30.00n
MM8 net120 net170 VDD VDD pch_mac W=120.00n L=30.00n
MM7 net186 cn net120 VDD pch_mac W=120.00n L=30.00n
MM5 net170 net186 VDD VDD pch_mac W=200.00n L=30.00n
MM15 net170 cn net161 VDD pch_mac W=0.2u L=30.00n
MM33 net186 c net126 VDD pch_mac W=0.2u L=30.00n
MM1 net126 D net129 VDD pch_mac W=200.00n L=30.00n
MM21 net146 net161 VDD VDD pch_mac W=200.00n L=30.00n
MM24 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM19 net89 net146 VDD VDD pch_mac W=120.00n L=30.00n
MM20 net161 c net89 VDD pch_mac W=120.00n L=30.00n
MM37 net137 SI VDD VDD pch_mac W=0.2u L=30.00n
MM36 net126 SEN net137 VDD pch_mac W=0.2u L=30.00n
MM31 net194 SI net198 VSS nch_mac W=0.2u L=30.00n
MM6 net186 c net162 VSS nch_mac W=120.00n L=30.00n
MM10 c CKN VSS VSS nch_mac W=0.2u L=30.00n
MM16 net154 net146 VSS VSS nch_mac W=120.00n L=30.00n
MM2 net190 D VSS VSS nch_mac W=200.00n L=30.00n
MM32 net186 cn net194 VSS nch_mac W=0.2u L=30.00n
MM25 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM30 net198 SE VSS VSS nch_mac W=0.2u L=30.00n
MM3 net194 SEN net190 VSS nch_mac W=200.00n L=30.00n
MM22 Q net146 VSS VSS nch_mac W=0.4u L=30.00n
MM18 net146 net161 VSS VSS nch_mac W=200.00n L=30.00n
MM17 net161 cn net154 VSS nch_mac W=120.00n L=30.00n
MM14 net170 c net161 VSS nch_mac W=0.2u L=30.00n
MM9 net162 net170 VSS VSS nch_mac W=120.00n L=30.00n
MM4 net170 net186 VSS VSS nch_mac W=0.2u L=30.00n
MM12 cn c VSS VSS nch_mac W=0.2u L=30.00n
.ENDS SNDQV4
.SUBCKT SNDRNQV4 CKN D Q RDN SE SI VDD VSS
MM34 SEN SE VDD VDD pch_mac W=0.2u L=30.00n
MM25 net107 RDN VDD VDD pch_mac W=0.2u L=30.00n
MM8 net107 net159 VDD VDD pch_mac W=120.00n L=30.00n
MM19 net98 net199 VDD VDD pch_mac W=120.00n L=30.00n
MM5 net159 net223 VDD VDD pch_mac W=200.00n L=30.00n
MM23 Q net199 VDD VDD pch_mac W=0.4u L=30.00n
MM7 net223 cn net107 VDD pch_mac W=0.2u L=30.00n
MM20 net198 c net98 VDD pch_mac W=120.00n L=30.00n
MM27 net199 RDN VDD VDD pch_mac W=200.00n L=30.00n
MM0 net150 SE VDD VDD pch_mac W=200.00n L=30.00n
MM36 net147 SEN net142 VDD pch_mac W=0.2u L=30.00n
MM37 net142 SI VDD VDD pch_mac W=0.2u L=30.00n
MM33 net223 c net147 VDD pch_mac W=0.2u L=30.00n
MM1 net147 D net150 VDD pch_mac W=200.00n L=30.00n
MM13 cn c VDD VDD pch_mac W=0.2u L=30.00n
MM15 net159 cn net198 VDD pch_mac W=0.2u L=30.00n
MM11 c CKN VDD VDD pch_mac W=200.00n L=30.00n
MM21 net199 net198 VDD VDD pch_mac W=200.00n L=30.00n
MM32 net223 cn net215 VSS nch_mac W=120.00n L=30.00n
MM31 net215 SI net211 VSS nch_mac W=0.2u L=30.00n
MM10 c CKN VSS VSS nch_mac W=0.2u L=30.00n
MM3 net215 SEN net219 VSS nch_mac W=200.00n L=30.00n
MM22 Q net199 VSS VSS nch_mac W=0.4u L=30.00n
MM6 net223 c net175 VSS nch_mac W=120.00n L=30.00n
MM18 net199 RDN net203 VSS nch_mac W=200.00n L=30.00n
MM16 net163 net199 VSS VSS nch_mac W=120.00n L=30.00n
MM30 net211 SE VSS VSS nch_mac W=0.2u L=30.00n
MM9 net175 net159 net179 VSS nch_mac W=120.00n L=30.00n
MM4 net159 net223 VSS VSS nch_mac W=0.2u L=30.00n
MM35 SEN SE VSS VSS nch_mac W=0.2u L=30.00n
MM17 net198 cn net163 VSS nch_mac W=120.00n L=30.00n
MM14 net159 c net198 VSS nch_mac W=0.2u L=30.00n
MM24 net179 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM12 cn c VSS VSS nch_mac W=0.2u L=30.00n
MM2 net219 D VSS VSS nch_mac W=200.00n L=30.00n
MM26 net203 net198 VSS VSS nch_mac W=200.00n L=30.00n
.ENDS SNDRNQV4
.SUBCKT SNDSRNQV4 CKN D Q RDN SDN SE SI VDD VSS
MM7 net106 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM8 net185 cn net106 VDD pch_mac W=120.00n L=30.00n
MM20 net189 c net166 VDD pch_mac W=120.00n L=30.00n
MM6 net106 net198 VDD VDD pch_mac W=120.00n L=30.00n
MM19 net166 net202 VDD VDD pch_mac W=120.00n L=30.00n
MM25 net166 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM40 SEN SE VDD VDD pch_mac W=120.00n L=30.00n
MM13 cn c VDD VDD pch_mac W=200.00n L=30.00n
MM11 c CKN VDD VDD pch_mac W=200.00n L=30.00n
MM23 Q net202 VDD VDD pch_mac W=400.00n L=30.00n
MM24 net198 SDN VDD VDD pch_mac W=120.00n L=30.00n
MM5 net198 net185 VDD VDD pch_mac W=200.00n L=30.00n
MM27 net202 RDN VDD VDD pch_mac W=120.00n L=30.00n
MM21 net202 net189 VDD VDD pch_mac W=200.00n L=30.00n
MM35 net190 SEN net133 VDD pch_mac W=120.00n L=30.00n
MM38 net190 D net129 VDD pch_mac W=200.00n L=30.00n
MM15 net198 cn net189 VDD pch_mac W=200.00n L=30.00n
MM0 net190 c net185 VDD pch_mac W=200.00n L=30.00n
MM36 net133 SI VDD VDD pch_mac W=120.00n L=30.00n
MM37 net129 SE VDD VDD pch_mac W=200.00n L=30.00n
MM14 net198 c net189 VSS nch_mac W=200.00n L=30.00n
MM3 net190 cn net185 VSS nch_mac W=200.00n L=30.00n
MM26 net226 SDN VSS VSS nch_mac W=200.00n L=30.00n
MM29 net178 SDN VSS VSS nch_mac W=120.00n L=30.00n
MM16 net174 net202 net178 VSS nch_mac W=120.00n L=30.00n
MM17 net189 cn net174 VSS nch_mac W=120.00n L=30.00n
MM18 net202 RDN net214 VSS nch_mac W=200.00n L=30.00n
MM2 net218 SI VSS VSS nch_mac W=120.00n L=30.00n
MM33 net210 SEN VSS VSS nch_mac W=200.00n L=30.00n
MM22 Q net202 VSS VSS nch_mac W=400.00n L=30.00n
MM1 net190 SE net218 VSS nch_mac W=120.00n L=30.00n
MM30 net214 net189 VSS VSS nch_mac W=200.00n L=30.00n
MM44 net222 RDN VSS VSS nch_mac W=120.00n L=30.00n
MM4 net198 net185 net226 VSS nch_mac W=200.00n L=30.00n
MM43 net230 net198 net222 VSS nch_mac W=120.00n L=30.00n
MM34 net190 D net210 VSS nch_mac W=200.00n L=30.00n
MM39 SEN SE VSS VSS nch_mac W=120.00n L=30.00n
MM9 net185 c net230 VSS nch_mac W=120.00n L=30.00n
MM12 cn c VSS VSS nch_mac W=200.00n L=30.00n
MM10 c CKN VSS VSS nch_mac W=200.00n L=30.00n
.ENDS SNDSRNQV4
.SUBCKT TBUFV4 I OE Z VDD VSS
MM43 net080 I VSS VSS nch_mac W=200.00n L=30.00n
MM44 net080 oen VSS VSS nch_mac W=200.00n L=30.00n
MM27 oen OE VSS VSS nch_mac W=120.00n L=30.00n
MM22 Z net080 VSS VSS nch_mac W=400.00n L=30.00n
MM36 net080 OE net_0163 VSS nch_mac W=200.00n L=30.00n
MM45 net_0163 OE VDD VDD pch_mac W=200.00n L=30.00n
MM46 net_0163 I VDD VDD pch_mac W=200.00n L=30.00n
MM28 oen OE VDD VDD pch_mac W=120.00n L=30.00n
MM21 Z net_0163 VDD VDD pch_mac W=400.00n L=30.00n
MM39 net080 oen net_0163 VDD pch_mac W=200.00n L=30.00n
.ENDS TBUFV4
.SUBCKT XNOR2V4 A1 A2 ZN VDD VSS
MM2 net30 A2 VDD VDD pch_mac W=200.00n L=30.00n
MM12 net29 A2 VDD VDD pch_mac W=400.00n L=30.00n
MM6 ZN net30 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net30 A1 VDD VDD pch_mac W=200.00n L=30.00n
MM13 ZN A1 net29 VDD pch_mac W=400.00n L=30.00n
MM16 net46 A1 VSS VSS nch_mac W=200.00n L=30.00n
MM15 net54 net30 VSS VSS nch_mac W=400.00n L=30.00n
MM8 ZN A1 net54 VSS nch_mac W=400.00n L=30.00n
MM14 ZN A2 net54 VSS nch_mac W=400.00n L=30.00n
MM17 net30 A2 net46 VSS nch_mac W=200.00n L=30.00n
.ENDS XNOR2V4
.SUBCKT XNOR3V4 A1 A2 A3 ZN VDD VSS
MMN1 net73 A1 VSS VSS nch_mac W=0.12u L=30.00n
MM19 net69 A2 VSS VSS nch_mac W=0.12u L=30.00n
MM16 net65 A3 VSS VSS nch_mac W=200.00n L=30.00n
MM22 net73 A2 VSS VSS nch_mac W=0.12u L=30.00n
MM20 MIDP net73 VSS VSS nch_mac W=0.12u L=30.00n
MM14 ZN MIDP net41 VSS nch_mac W=400.000n L=30.00n
MM15 net41 net120 VSS VSS nch_mac W=400.000n L=30.00n
MM17 net120 MIDP net65 VSS nch_mac W=200.00n L=30.00n
MM11 MIDP A1 net69 VSS nch_mac W=0.12u L=30.00n
MM8 ZN A3 net41 VSS nch_mac W=400.000n L=30.00n
MM12 net88 MIDP VDD VDD pch_mac W=400.00n L=30.00n
MM6 ZN net120 VDD VDD pch_mac W=400.00n L=30.00n
MM5 net120 MIDP VDD VDD pch_mac W=200.00n L=30.00n
MM9 net73 A2 net80 VDD pch_mac W=0.12u L=30.00n
MM0 MIDP A1 net96 VDD pch_mac W=0.145u L=30.00n
MM13 ZN A3 net88 VDD pch_mac W=400.00n L=30.00n
MM2 net120 A3 VDD VDD pch_mac W=200.00n L=30.00n
MM10 net80 A1 VDD VDD pch_mac W=0.12u L=30.00n
MM1 MIDP A2 net96 VDD pch_mac W=0.145u L=30.00n
MM3 net96 net73 VDD VDD pch_mac W=0.12u L=30.00n
.ENDS XNOR3V4
.SUBCKT XOR2V4 A1 A2 Z VDD VSS
MMN1 net39 A1 VSS VSS nch_mac W=200.00n L=30.00n
MM1 net39 A2 VSS VSS nch_mac W=200.00n L=30.00n
MM0 Z A1 net27 VSS nch_mac W=400.00n L=30.00n
MM5 net27 A2 VSS VSS nch_mac W=400.00n L=30.00n
MM2 Z net39 VSS VSS nch_mac W=400.00n L=30.00n
MM12 net58 net39 VDD VDD pch_mac W=400.00n L=30.00n
MM13 Z A2 net58 VDD pch_mac W=400.00n L=30.00n
MM3 net46 A1 VDD VDD pch_mac W=200.00n L=30.00n
MM6 Z A1 net58 VDD pch_mac W=400.00n L=30.00n
MM8 net39 A2 net46 VDD pch_mac W=200.00n L=30.00n
.ENDS XOR2V4
.SUBCKT XOR3V4 A1 A2 A3 Z VDD VSS
MM11 net52 A1 VDD VDD pch_mac W=0.12u L=30.00n
MM26 Z net36 VDD VDD pch_mac W=400.00n L=30.00n
MM24 net75 MIDP VDD VDD pch_mac W=400.00n L=30.00n
MM23 net36 A3 VDD VDD pch_mac W=200.00n L=30.00n
MM22 net36 MIDP VDD VDD pch_mac W=200.00n L=30.00n
MM25 Z A3 net75 VDD pch_mac W=400.00n L=30.00n
MM4 net52 A2 VDD VDD pch_mac W=0.12u L=30.00n
MM12 net63 A2 VDD VDD pch_mac W=0.12u L=30.00n
MM13 MIDP A1 net63 VDD pch_mac W=0.12u L=30.00n
MM6 MIDP net52 VDD VDD pch_mac W=0.12u L=30.00n
MM20 Z MIDP net108 VSS nch_mac W=400.000n L=30.00n
MM19 net108 net36 VSS VSS nch_mac W=400.000n L=30.00n
MM21 Z A3 net108 VSS nch_mac W=400.000n L=30.00n
MM15 net36 MIDP net92 VSS nch_mac W=200.00n L=30.00n
MMN1 net96 A1 VSS VSS nch_mac W=0.12u L=30.00n
MM16 net92 A3 VSS VSS nch_mac W=200.00n L=30.00n
MM9 MIDP A2 net84 VSS nch_mac W=0.145u L=30.00n
MM7 net84 net52 VSS VSS nch_mac W=0.12u L=30.00n
MM5 MIDP A1 net84 VSS nch_mac W=0.145u L=30.00n
MM14 net52 A2 net96 VSS nch_mac W=0.12u L=30.00n
.ENDS XOR3V4
